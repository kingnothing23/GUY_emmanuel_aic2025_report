* NGSPICE file created from JNW_GR01.ext - technology: sky130A

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt JNW_GR01 VDD vref cmp reset VSS
*.subckt JNW_GR01 VDD VSS reset cmp vref
X0 VDD xa1.xe1.G xa1.xb1.S VDD sky130_fd_pr__pfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X1 VDD xb1.xa2.P cmp VDD sky130_fd_pr__pfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X2 a_14460_6992# a_14676_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X3 xa1.xa2.xc1.D xa1.xb1.S xa1.xa2.xc2.G VSS sky130_fd_pr__nfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X4 xb1.xb3.G vref xb1.xb2.S xb1.xb2.S sky130_fd_pr__pfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X5 VSS xb1.xb3.D cmp VSS sky130_fd_pr__nfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X6 VDD xa1.xa2.xd1.D xa1.xe1.G VDD sky130_fd_pr__pfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X7 xa1.xa2.xc1.D xa1.xa2.xa1.G VSS VSS sky130_fd_pr__nfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X8 VSS xb1.xb3.G xb1.xb3.G VSS sky130_fd_pr__nfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X9 xa1.xa2.xa1.G xa1.xa2.xa1.G VSS VSS sky130_fd_pr__nfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X10 cmp xb1.xe.D sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X11 vref xa1.xe1.G VDD VDD sky130_fd_pr__pfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X12 VDD xa1.xe1.G xb3.A VDD sky130_fd_pr__pfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X13 VSS VSS xa1.xb1.S VDD sky130_fd_pr__pfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X14 VSS xa1.xe1.G sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X15 VSS xa1.xe1.G sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X16 cmp xb1.xa2.P VDD VDD sky130_fd_pr__pfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
X17 a_1660_3480# a_1876_1560# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X18 VDD xa1.xa2.xc2.G xa1.xa2.xd1.D VDD sky130_fd_pr__pfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X19 xb1.xb3.G xb1.xb3.G VSS VSS sky130_fd_pr__nfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
X20 cmp xb1.xb3.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
X21 xa1.xb1.S xa1.xe1.G VDD VDD sky130_fd_pr__pfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X22 a_10580_5712# a_10364_3792# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X23 a_15756_6992# a_15972_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X24 a_16188_6992# a_15972_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X25 xb3.A reset VSS VSS sky130_fd_pr__nfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X26 a_10148_5712# a_10364_3792# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X27 a_796_3480# a_580_1560# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X28 a_15756_6992# a_15540_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X29 VDD xa1.xa2.xc2.G xa1.xa2.xc2.G VDD sky130_fd_pr__pfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X30 VSS xa1.xa2.xa1.G xa1.xe1.G VSS sky130_fd_pr__nfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X31 a_10148_5712# a_9932_3792# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X32 a_14460_6992# a_14244_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X33 xb1.xb3.D xb1.xb3.G VSS VSS sky130_fd_pr__nfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
X34 VDD xb1.xa2.P xb1.xa2.P VDD sky130_fd_pr__pfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X35 VSS xa1.xe1.G sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X36 VSS xa1.xe1.G sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X37 VSS VSS xa1.xb2.S VDD sky130_fd_pr__pfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X38 VSS a_14244_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X39 xa1.xa2.xd1.D xa1.xc1.P xa1.xa2.xc1.D VSS sky130_fd_pr__nfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X40 xa1.xb2.S a_9500_280# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X41 xb1.xb3.D xb3.A xb1.xb2.S xb1.xb2.S sky130_fd_pr__pfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X42 VDD a_1876_1560# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X43 xb1.xa2.N a_17268_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X44 xb1.xa2.P xb1.xa2.P VDD VDD sky130_fd_pr__pfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
X45 xb1.xb2.S vref xb1.xb3.G xb1.xb2.S sky130_fd_pr__pfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X46 xb1.xb3.D VDD xb1.xe.D VSS sky130_fd_pr__nfet_01v8 ad=0.4704 pd=2.9 as=0.2784 ps=1.54 w=0.96 l=0.22
X47 a_1660_3480# a_1444_1560# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X48 a_9716_5712# a_9932_3792# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X49 a_17052_6992# a_17268_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X50 VSS xa1.xa2.xa1.G xa1.xa2.xc1.D VSS sky130_fd_pr__nfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X51 VDD xa1.xe1.G vref VDD sky130_fd_pr__pfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X52 a_16620_6992# a_16836_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X53 VSS xa1.xa2.xa1.G xa1.xa2.xa1.G VSS sky130_fd_pr__nfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X54 xa1.xe1.G xa1.xa2.xd1.D VDD VDD sky130_fd_pr__pfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X55 a_1228_3480# a_1444_1560# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X56 a_9716_5712# a_9500_3792# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X57 VDD xb1.xa2.P xb1.xb2.S VDD sky130_fd_pr__pfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X58 xa1.xa2.xa1.G a_580_1560# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X59 a_1228_3480# a_1012_1560# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X60 a_15324_6992# a_15540_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X61 xa1.xb1.S VSS VSS VDD sky130_fd_pr__pfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X62 xb1.xa2.P a_14244_1560# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X63 xa1.xc1.P a_9500_280# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X64 xb3.A xa1.xe1.G VDD VDD sky130_fd_pr__pfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X65 xb1.xe.D VDD xb1.xb3.D VSS sky130_fd_pr__nfet_01v8 ad=0.2784 pd=1.54 as=0.4704 ps=2.9 w=0.96 l=0.22
X66 a_15324_6992# a_15108_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X67 xb1.xa2.N a_14244_1560# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X68 VSS reset xb3.A VSS sky130_fd_pr__nfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X69 a_14892_6992# a_15108_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X70 xa1.xa2.xd1.D xa1.xa2.xc2.G VDD VDD sky130_fd_pr__pfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X71 xa1.xa2.xc2.G xa1.xb1.S xa1.xa2.xc1.D VSS sky130_fd_pr__nfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X72 VSS xb3.A sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X73 a_17052_6992# a_16836_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X74 xa1.xa2.xc2.G xa1.xa2.xc2.G VDD VDD sky130_fd_pr__pfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X75 xa1.xb2.S VSS VSS VDD sky130_fd_pr__pfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X76 xa1.xa2.xc1.D xa1.xc1.P xa1.xa2.xd1.D VSS sky130_fd_pr__nfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X77 a_16620_6992# a_16404_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X78 xa1.xe1.G xa1.xa2.xa1.G VSS VSS sky130_fd_pr__nfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X79 xa1.xc1.P a_9500_3792# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X80 a_10580_5712# a_10796_3792# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X81 xb1.xb2.S xb3.A xb1.xb3.D xb1.xb2.S sky130_fd_pr__pfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X82 vref a_10796_3792# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X83 a_16188_6992# a_16404_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X84 VSS xb1.xb3.G xb1.xb3.D VSS sky130_fd_pr__nfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X85 xa1.xe1.G xa1.xa2.xd1.D sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X86 a_796_3480# a_1012_1560# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X87 a_14892_6992# a_14676_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X88 xb1.xb2.S xb1.xa2.P VDD VDD sky130_fd_pr__pfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
C0 a_15656_9378# xb1.xe.D 0.02838f
C1 xa1.xb1.S a_7248_1258# 0.05989f
C2 a_160_11138# vref 0.01375f
C3 xa1.xa2.xc1.D xa1.xa2.xa1.G 0.39846f
C4 xb1.xa2.N xb3.A 0.08653f
C5 a_18976_1258# xb3.A 0.07043f
C6 a_14460_6992# a_14892_6992# 0.21349f
C7 a_18976_2320# a_18976_2480# 0.11476f
C8 xa1.xa2.xd1.D xa1.xe1.G 3.66269f
C9 a_18976_586# a_18976_746# 0.11476f
C10 a_14244_5072# a_14028_5072# 0.01515f
C11 xa1.xa2.xc1.D a_3584_1000# 0.03962f
C12 xa1.xa2.xc1.D xa1.xb1.S 0.62862f
C13 xb3.A a_18976_2058# 0.07261f
C14 a_13824_9858# a_13824_10018# 0.11476f
C15 a_3584_3114# xa1.xb1.S 0.07921f
C16 xa1.xa2.xc2.G xa1.xa2.xa1.G 0.06798f
C17 a_3480_7164# VDD 0.04426f
C18 xa1.xa2.xa1.G a_3584_200# 0.07059f
C19 a_11228_3792# a_10796_3792# 0.01515f
C20 cmp a_13824_10018# 0.02114f
C21 xb1.xa2.P a_15756_6992# 0.12598f
C22 xb1.xb2.S a_18976_106# 0.03384f
C23 xa1.xc1.P a_5416_188# 0.07046f
C24 a_13824_944# xb1.xa2.P 0.11958f
C25 xa1.xa2.xc2.G xa1.xb1.S 0.44796f
C26 cmp a_13824_9218# 0.01491f
C27 xb1.xb2.S xb1.xb3.G 0.78799f
C28 a_14028_5072# xb1.xa2.N 0.10537f
C29 VDD a_14676_5072# 0.0263f
C30 a_15656_9218# xb1.xb3.D 0.02923f
C31 xb1.xb3.D a_15756_6992# 0.01142f
C32 a_13824_11898# a_13824_12378# 0.03053f
C33 cmp xb1.xe.D 3.29556f
C34 reset xb1.xb3.D 0.03025f
C35 xb1.xb3.D xb1.xa2.P 0.02783f
C36 xa1.xa2.xa1.G a_3584_1000# 0.07255f
C37 xa1.xb1.S xa1.xa2.xa1.G 0.19245f
C38 xb1.xe.D a_15656_10018# 0.02333f
C39 a_16404_5072# a_15972_5072# 0.14233f
C40 xa1.xc1.P a_9932_280# 0.02416f
C41 xa1.xc1.P xa1.xa2.xc1.D 1.05094f
C42 a_15656_9858# xb1.xe.D 0.02992f
C43 xb1.xa2.N a_17700_5072# 0.1466f
C44 xb1.xa2.N xb1.xa2.P 0.58692f
C45 a_15656_9378# VDD 0.08135f
C46 VDD a_14892_6992# 0.01333f
C47 VDD a_3584_2058# 0.48562f
C48 xa1.xa2.xd1.D a_5416_988# 0.03482f
C49 a_14676_1560# a_14244_1560# 0.01515f
C50 a_13824_11738# xb1.xb3.D 0.08445f
C51 a_11228_3792# VDD 0.0154f
C52 a_14244_5072# xb1.xa2.N 0.21356f
C53 xa1.xa2.xc2.G xa1.xc1.P 0.29273f
C54 a_160_9538# VDD 0.63332f
C55 a_10580_5712# a_10148_5712# 0.21349f
C56 xb3.A a_13824_12378# 0.01825f
C57 VDD a_3584_2314# 0.05433f
C58 xb1.xa2.N xb1.xb3.D 0.02365f
C59 a_18976_1258# xb1.xb3.D 0.013f
C60 a_13824_11098# a_13824_10018# 0.01285f
C61 xb1.xb2.S vref 3.32417f
C62 a_364_1560# a_580_1560# 0.01515f
C63 a_1228_3480# a_796_3480# 0.21349f
C64 xb1.xe.D vref 0.13557f
C65 xb1.xb2.S a_20808_1514# 0.05316f
C66 a_1012_1560# a_580_1560# 0.14233f
C67 a_160_11138# xb3.A 0.01377f
C68 a_18976_2058# xb1.xb3.D 0.03695f
C69 a_3480_8232# VDD 0.63595f
C70 a_18976_3120# xb1.xb3.D 0.02778f
C71 a_14460_6992# vref 0.01128f
C72 a_18976_106# VDD 0.50265f
C73 xa1.xc1.P xa1.xa2.xa1.G 0.0186f
C74 xa1.xb1.S a_7248_458# 0.05903f
C75 xa1.xc1.P a_9716_5712# 0.24739f
C76 a_10580_5712# VDD 0.08469f
C77 a_5416_1258# VDD 0.4831f
C78 a_18976_2320# xb1.xb3.G 0.02601f
C79 a_13824_11098# xb1.xe.D 0.02468f
C80 a_18976_1258# a_18976_746# 0.02844f
C81 a_20808_2154# xb1.xb3.G 0.11839f
C82 xa1.xc1.P xa1.xb1.S 0.31142f
C83 VDD a_13824_9858# 0.49339f
C84 xa1.xa2.xd1.D a_5416_188# 0.013f
C85 cmp VDD 1.01572f
C86 a_14676_1560# xb1.xa2.P 0.245f
C87 xb1.xb3.G a_18976_2480# 0.08513f
C88 a_3480_7432# VDD 0.48236f
C89 a_15972_5072# xb1.xa2.P 0.01443f
C90 VDD a_15656_9858# 0.08122f
C91 xa1.xa2.xc2.G a_5416_2058# 0.07197f
C92 a_3584_1258# xa1.xa2.xc1.D 0.02378f
C93 a_13824_9378# a_13824_9218# 0.11476f
C94 a_9284_3792# xa1.xc1.P 0.16915f
C95 reset a_13824_12378# 0.07043f
C96 a_3480_7164# a_3480_7432# 0.05943f
C97 xa1.xa2.xd1.D xa1.xa2.xc1.D 0.40891f
C98 VDD xa1.xe1.G 8.65756f
C99 a_3480_6364# xa1.xe1.G 0.016f
C100 a_14028_1560# a_14244_1560# 0.01515f
C101 a_13824_464# VDD 0.50552f
C102 a_20808_1674# a_20808_2154# 0.01174f
C103 xa1.xa2.xc2.G a_3584_1258# 0.08851f
C104 a_3584_2314# a_3584_2058# 0.06279f
C105 a_20808_458# xb1.xb2.S 0.6232f
C106 a_15108_5072# xb1.xa2.P 0.02072f
C107 VDD vref 3.11495f
C108 xa1.xa2.xc2.G xa1.xa2.xd1.D 0.37323f
C109 a_18976_2960# a_18976_2480# 0.01174f
C110 xb1.xb3.D a_13824_12378# 0.01721f
C111 xb1.xa2.P a_15540_5072# 0.30811f
C112 a_3480_7164# xa1.xe1.G 0.07424f
C113 xb1.xa2.N a_15972_5072# 0.02767f
C114 a_7248_1258# xa1.xb2.S 0.05639f
C115 a_160_1160# xa1.xa2.xa1.G 0.09668f
C116 a_364_1560# xa1.xa2.xa1.G 0.05799f
C117 a_9284_280# xa1.xb2.S 0.01797f
C118 xb1.xb2.S a_18976_586# 0.03571f
C119 a_1012_1560# xa1.xa2.xa1.G 0.03175f
C120 xb1.xb2.S xb3.A 2.5859f
C121 a_3584_1258# a_3584_1000# 0.06221f
C122 a_16188_6992# vref 0.01128f
C123 xa1.xa2.xd1.D xa1.xa2.xa1.G 0.66101f
C124 xb3.A xb1.xe.D 0.01028f
C125 a_1660_3480# VDD 0.21862f
C126 a_1876_1560# a_2308_1560# 0.01515f
C127 xa1.xa2.xa1.G a_796_3480# 0.30226f
C128 a_14028_1560# xb1.xa2.P 0.04127f
C129 xa1.xa2.xd1.D xa1.xb1.S 0.49431f
C130 a_16620_6992# a_16188_6992# 0.21349f
C131 xb1.xa2.N a_15108_5072# 0.03028f
C132 cmp a_13824_11258# 0.0414f
C133 xb1.xa2.N a_15540_5072# 0.0171f
C134 a_9284_280# a_9500_280# 0.01515f
C135 a_9500_280# a_9932_280# 0.01515f
C136 a_160_10338# VDD 0.59061f
C137 xb1.xb2.S a_20808_1258# 0.4835f
C138 VDD a_5416_988# 0.04502f
C139 a_160_11938# VDD 0.62226f
C140 VDD a_13824_9378# 0.50229f
C141 a_160_9538# xa1.xe1.G 0.08355f
C142 cmp a_13824_9858# 0.03718f
C143 xa1.xb1.S xa1.xb2.S 0.19242f
C144 a_14892_6992# vref 0.01128f
C145 a_14028_1560# xb1.xa2.N 0.01537f
C146 a_13824_9218# xb1.xa2.P 0.02164f
C147 a_11228_3792# vref 0.01683f
C148 a_15656_9218# xb1.xe.D 0.01169f
C149 a_17268_5072# a_16836_5072# 0.14233f
C150 a_13824_304# VDD 0.58305f
C151 xb1.xb2.S xb1.xa2.P 0.18817f
C152 xa1.xa2.xd1.D xa1.xc1.P 0.46738f
C153 a_3480_8232# xa1.xe1.G 0.01492f
C154 xb1.xe.D xb1.xa2.P 0.03409f
C155 a_1444_1560# xa1.xa2.xa1.G 0.01378f
C156 a_18976_586# VDD 0.49275f
C157 a_2308_1560# VDD 0.02278f
C158 a_15656_9858# a_15656_10018# 0.0971f
C159 xb3.A VDD 0.97855f
C160 a_15324_6992# a_14892_6992# 0.21349f
C161 a_1876_1560# xa1.xa2.xa1.G 0.01584f
C162 xb1.xb3.G a_18976_2960# 0.08185f
C163 a_13824_11098# a_13824_11258# 0.11476f
C164 xb1.xb2.S xb1.xb3.D 0.82144f
C165 a_13824_1104# xb1.xa2.P 0.07112f
C166 a_13824_944# a_13824_1104# 0.11476f
C167 a_20808_1674# xb1.xb3.G 0.11472f
C168 a_10580_5712# vref 0.23257f
C169 xb1.xb3.D xb1.xe.D 0.78734f
C170 a_15972_5072# a_15540_5072# 0.14233f
C171 VDD a_7248_1258# 0.46453f
C172 VDD a_14244_1560# 0.06277f
C173 xb1.xb3.G vref 0.56812f
C174 a_3480_7432# xa1.xe1.G 0.06791f
C175 xa1.xc1.P xa1.xb2.S 0.3747f
C176 cmp vref 0.08918f
C177 xb1.xb2.S a_18976_1258# 0.50479f
C178 xb1.xb3.G a_20808_1514# 0.03885f
C179 a_9284_280# VDD 0.02515f
C180 a_14028_1560# a_14676_1560# 0.06667f
C181 xa1.xa2.xc1.D VDD 0.70229f
C182 xb1.xb2.S a_18976_746# 0.03533f
C183 a_14028_5072# VDD 0.09304f
C184 xb1.xb2.S a_18976_2058# 0.48226f
C185 cmp a_13824_11098# 0.08197f
C186 a_15108_5072# a_15540_5072# 0.14233f
C187 xa1.xa2.xc2.G VDD 6.13956f
C188 xa1.xa2.xd1.D a_5416_2058# 0.0376f
C189 a_10148_5712# a_9716_5712# 0.21349f
C190 a_9284_3792# a_9500_3792# 0.01515f
C191 a_15656_9218# VDD 0.01578f
C192 xa1.xe1.G vref 0.45178f
C193 a_5416_1258# a_5416_988# 0.0589f
C194 VDD xb1.xa2.P 8.73304f
C195 a_13824_944# VDD 0.50687f
C196 a_20808_1674# a_20808_1514# 0.11476f
C197 VDD xa1.xa2.xa1.G 0.32684f
C198 xa1.xa2.xa1.G a_3480_6364# 0.08127f
C199 VDD a_9716_5712# 0.08362f
C200 xa1.xc1.P a_9500_3792# 0.14826f
C201 a_14244_5072# VDD 0.03646f
C202 a_18976_2320# xb1.xb3.D 0.03393f
C203 xa1.xc1.P a_9932_3792# 0.19092f
C204 VDD a_3584_1000# 0.05123f
C205 a_16188_6992# a_15756_6992# 0.21349f
C206 a_13824_9378# a_13824_9858# 0.01174f
C207 xa1.xb1.S VDD 5.52295f
C208 cmp a_13824_11898# 0.01307f
C209 a_17268_5072# xb3.A 0.01159f
C210 VDD xb1.xb3.D 0.56002f
C211 a_16620_6992# vref 0.01128f
C212 cmp a_13824_9378# 0.03221f
C213 a_3480_7164# xa1.xa2.xa1.G 0.07043f
C214 a_20808_458# xb1.xb3.G 0.013f
C215 xb1.xb3.D a_18976_2480# 0.03329f
C216 a_15324_6992# vref 0.01067f
C217 a_18976_106# a_18976_586# 0.01174f
C218 xb1.xa2.N VDD 0.93258f
C219 a_18976_1258# VDD 0.02387f
C220 xa1.xa2.xc1.D a_3584_2058# 0.01931f
C221 a_16188_6992# xb1.xb3.D 0.01324f
C222 a_160_10338# xa1.xe1.G 0.14277f
C223 a_18976_2320# a_18976_2058# 0.06106f
C224 VDD a_18976_746# 0.42427f
C225 a_14244_5072# a_14676_5072# 0.14233f
C226 a_160_11938# xa1.xe1.G 0.07043f
C227 xb1.xb3.G xb3.A 0.0992f
C228 xa1.xa2.xc1.D a_3584_2314# 0.07083f
C229 VDD a_7248_458# 0.56587f
C230 xa1.xa2.xc2.G a_3584_2058# 0.12259f
C231 a_160_10338# vref 0.01571f
C232 cmp xb3.A 0.63749f
C233 a_15656_9218# a_15656_9378# 0.0971f
C234 xa1.xc1.P VDD 1.11748f
C235 xa1.xa2.xc2.G a_3584_2314# 0.04553f
C236 a_14892_6992# xb1.xa2.P 0.01614f
C237 a_5416_1258# xa1.xa2.xc1.D 0.0142f
C238 xb3.A a_13824_13178# 0.05579f
C239 a_1444_1560# a_1012_1560# 0.14233f
C240 a_17052_6992# vref 0.01128f
C241 a_20808_2154# a_20808_2314# 0.11476f
C242 xb1.xa2.N a_14676_5072# 0.03684f
C243 a_13824_304# a_13824_464# 0.11476f
C244 a_17268_5072# a_17700_5072# 0.01515f
C245 a_20808_1258# xb1.xb3.G 0.03814f
C246 a_20808_458# vref 0.09933f
C247 xb1.xb2.S a_18976_n54# 0.01206f
C248 xb3.A xa1.xe1.G 0.44469f
C249 a_15656_9378# xb1.xb3.D 0.05643f
C250 xa1.xa2.xc2.G a_5416_1258# 0.07046f
C251 a_14676_1560# VDD 0.04628f
C252 a_16620_6992# a_17052_6992# 0.21349f
C253 a_16404_5072# a_16836_5072# 0.14233f
C254 a_1660_3480# a_1228_3480# 0.21349f
C255 a_160_9538# xa1.xb1.S 0.03503f
C256 a_18976_106# xb1.xa2.P 0.08182f
C257 a_13824_11258# xb1.xb3.D 0.08168f
C258 xb3.A vref 1.53064f
C259 xa1.xb1.S a_3584_2314# 0.07117f
C260 a_13824_11738# a_13824_11258# 0.01174f
C261 a_7248_2058# xa1.xb2.S 0.08238f
C262 xb1.xa2.P a_13824_9858# 0.08107f
C263 reset cmp 0.08768f
C264 a_17268_5072# xb1.xa2.N 0.02892f
C265 cmp xb1.xa2.P 0.22101f
C266 VDD a_5416_2058# 0.63014f
C267 xb1.xe.D a_13824_10018# 0.03353f
C268 a_160_11138# VDD 0.58707f
C269 a_20808_1258# vref 0.07201f
C270 xb1.xb3.G xb1.xb3.D 0.43731f
C271 reset a_13824_13178# 0.07043f
C272 VDD a_15108_5072# 0.01168f
C273 cmp xb1.xb3.D 0.41757f
C274 a_20808_1258# a_20808_1514# 0.06279f
C275 a_3584_1258# VDD 0.48244f
C276 cmp a_13824_11738# 0.0349f
C277 xb1.xb3.D a_15656_10018# 0.0371f
C278 xa1.xa2.xd1.D VDD 4.24367f
C279 a_1876_1560# a_1444_1560# 0.14233f
C280 xa1.xa2.xd1.D a_3480_6364# 0.03942f
C281 a_15656_9858# xb1.xb3.D 0.05554f
C282 a_13824_464# xb1.xa2.P 0.11964f
C283 a_13824_464# a_13824_944# 0.01174f
C284 xa1.xa2.xa1.G xa1.xe1.G 0.49041f
C285 a_18976_n54# VDD 0.58137f
C286 a_15756_6992# vref 0.01128f
C287 a_160_11938# xb3.A 0.0156f
C288 xb1.xb3.G a_18976_2058# 0.01323f
C289 xb1.xa2.P vref 0.237f
C290 xa1.xb1.S xa1.xe1.G 0.49818f
C291 a_14028_1560# VDD 0.0554f
C292 a_17052_6992# xb3.A 0.012f
C293 a_18976_2960# xb1.xb3.D 0.02933f
C294 a_3480_7164# xa1.xa2.xd1.D 0.01088f
C295 a_15108_5072# a_14676_5072# 0.14233f
C296 xa1.xa2.xc1.D a_5416_988# 0.08009f
C297 xa1.xb1.S vref 0.08264f
C298 xb1.xb3.D vref 1.41264f
C299 a_9932_3792# a_9500_3792# 0.14233f
C300 VDD xa1.xb2.S 0.92687f
C301 a_10796_3792# a_10364_3792# 0.14233f
C302 a_15324_6992# a_15756_6992# 0.21349f
C303 xb1.xb3.G a_20808_2314# 0.05596f
C304 a_10364_3792# a_9932_3792# 0.14233f
C305 xa1.xa2.xa1.G a_160_360# 0.1391f
C306 a_15324_6992# xb1.xa2.P 0.23404f
C307 a_1660_3480# xa1.xa2.xa1.G 0.01519f
C308 VDD a_13824_10018# 0.40658f
C309 a_16620_6992# xb1.xb3.D 0.01324f
C310 xb1.xa2.N a_16836_5072# 0.02767f
C311 xb1.xa2.N vref 0.01533f
C312 a_18976_3120# a_18976_2960# 0.11476f
C313 VDD a_13824_9218# 0.56296f
C314 xb1.xb2.S a_18976_2320# 0.04804f
C315 VDD a_7248_2058# 0.56635f
C316 xb1.xb2.S VDD 1.16666f
C317 VDD xb1.xe.D 0.44006f
C318 xa1.xa2.xc1.D a_5416_188# 0.0565f
C319 a_13824_9378# xb1.xa2.P 0.08242f
C320 a_14460_6992# VDD 0.0269f
C321 xa1.xc1.P vref 0.02744f
C322 xa1.xb1.S a_160_10338# 0.01299f
C323 xa1.xa2.xa1.G a_1228_3480# 0.02131f
C324 a_13824_1104# VDD 0.41828f
C325 a_13824_11898# xb1.xb3.D 0.0288f
C326 xa1.xa2.xa1.G a_580_1560# 0.10652f
C327 a_13824_304# xb1.xa2.P 0.05442f
C328 a_13824_11738# a_13824_11898# 0.11476f
C329 xa1.xa2.xd1.D a_3480_8232# 0.0713f
C330 a_9284_280# a_9932_280# 0.06667f
C331 a_17052_6992# xb1.xb3.D 0.01324f
C332 a_18976_586# xb1.xa2.P 0.08074f
C333 xa1.xa2.xd1.D a_5416_1258# 0.03715f
C334 reset xb3.A 0.77478f
C335 a_18976_n54# a_18976_106# 0.11476f
C336 xb3.A a_17700_5072# 0.01373f
C337 xa1.xa2.xc1.D a_3584_3114# 0.05775f
C338 a_2308_1560# xa1.xa2.xa1.G 0.03096f
C339 xb1.xa2.N a_17052_6992# 0.2491f
C340 a_10148_5712# VDD 0.08362f
C341 xa1.xa2.xc2.G xa1.xa2.xc1.D 1.38183f
C342 a_2308_1560# xa1.xb1.S 0.01722f
C343 xa1.xa2.xc1.D a_3584_200# 0.01326f
C344 xa1.xa2.xc2.G a_3584_3114# 0.01512f
C345 a_14244_1560# xb1.xa2.P 0.22449f
C346 xa1.xc1.P a_5416_988# 0.07237f
C347 a_160_11138# xa1.xe1.G 0.14277f
C348 xb3.A xb1.xb3.D 0.655f
C349 xa1.xa2.xd1.D a_3480_7432# 0.08395f
C350 a_16404_5072# xb1.xa2.N 0.02767f
C351 cmp VSS 9.49424f
C352 vref VSS 26.0141f
C353 reset VSS 5.2369f
C354 VDD VSS 0.1055p
C355 a_20808_458# VSS 0.02653f $ **FLOATING
C356 a_18976_n54# VSS 0.02916f $ **FLOATING
C357 a_18976_746# VSS 0.07212f $ **FLOATING
C358 a_13824_304# VSS 0.02981f $ **FLOATING
C359 a_20808_1258# VSS 0.05294f $ **FLOATING
C360 a_13824_1104# VSS 0.13937f $ **FLOATING
C361 a_18976_1258# VSS 0.07213f $ **FLOATING
C362 a_20808_1514# VSS 0.41005f $ **FLOATING
C363 a_20808_1674# VSS 0.49626f $ **FLOATING
C364 a_18976_2058# VSS 0.05665f $ **FLOATING
C365 a_20808_2154# VSS 0.50871f $ **FLOATING
C366 a_20808_2314# VSS 0.61822f $ **FLOATING
C367 a_18976_2320# VSS 0.41618f $ **FLOATING
C368 a_18976_2480# VSS 0.49887f $ **FLOATING
C369 xb1.xb3.G VSS 5.44947f
C370 a_18976_2960# VSS 0.50822f $ **FLOATING
C371 a_18976_3120# VSS 0.60866f $ **FLOATING
C372 a_14676_1560# VSS 1.82365f $ **FLOATING
C373 a_14244_1560# VSS 0.62373f
C374 a_14028_1560# VSS 1.83048f $ **FLOATING
C375 a_9932_280# VSS 1.86269f $ **FLOATING
C376 a_9500_280# VSS 0.6339f
C377 a_9284_280# VSS 1.82457f $ **FLOATING
C378 a_7248_458# VSS 0.15377f $ **FLOATING
C379 a_5416_188# VSS 0.58441f $ **FLOATING
C380 a_5416_988# VSS 0.4362f $ **FLOATING
C381 a_3584_200# VSS 0.67275f $ **FLOATING
C382 a_3584_1000# VSS 0.49132f $ **FLOATING
C383 a_160_360# VSS 0.6245f $ **FLOATING
C384 a_7248_1258# VSS 0.18787f $ **FLOATING
C385 a_160_1160# VSS 0.67829f $ **FLOATING
C386 xa1.xb2.S VSS 2.79865f
C387 a_7248_2058# VSS 0.10925f $ **FLOATING
C388 a_5416_1258# VSS 0.05098f $ **FLOATING
C389 a_5416_2058# VSS 0.02527f $ **FLOATING
C390 a_3584_1258# VSS 0.05879f $ **FLOATING
C391 a_3584_2058# VSS 0.04789f $ **FLOATING
C392 a_3584_2314# VSS 0.42696f $ **FLOATING
C393 xa1.xa2.xc2.G VSS 1.35097f
C394 xa1.xa2.xc1.D VSS 1.69501f
C395 a_3584_3114# VSS 0.58654f $ **FLOATING
C396 a_17700_5072# VSS 1.99287f $ **FLOATING
C397 xb1.xa2.N VSS 5.02623f
C398 a_17268_5072# VSS 0.5397f
C399 a_17052_6992# VSS 0.64011f
C400 a_16836_5072# VSS 0.44449f
C401 a_16620_6992# VSS 0.63998f
C402 a_16404_5072# VSS 0.44331f
C403 a_16188_6992# VSS 0.63914f
C404 a_15972_5072# VSS 0.44299f
C405 a_15756_6992# VSS 0.6436f
C406 a_15540_5072# VSS 0.43952f
C407 a_15324_6992# VSS 0.64723f
C408 a_15108_5072# VSS 0.44559f
C409 a_14892_6992# VSS 0.66546f
C410 a_14676_5072# VSS 0.44301f
C411 a_14460_6992# VSS 0.91526f
C412 a_14244_5072# VSS 0.53659f
C413 a_14028_5072# VSS 2.02206f $ **FLOATING
C414 a_11228_3792# VSS 1.91966f $ **FLOATING
C415 a_10796_3792# VSS 0.53218f
C416 a_10580_5712# VSS 0.63706f
C417 a_10364_3792# VSS 0.44635f
C418 a_10148_5712# VSS 0.63197f
C419 a_9932_3792# VSS 0.43595f
C420 a_9716_5712# VSS 0.63171f
C421 a_9500_3792# VSS 0.52984f
C422 xa1.xc1.P VSS 8.73835f
C423 a_9284_3792# VSS 1.89226f $ **FLOATING
C424 a_2308_1560# VSS 1.91857f $ **FLOATING
C425 a_1876_1560# VSS 0.54859f
C426 a_1660_3480# VSS 0.64331f
C427 a_1444_1560# VSS 0.45225f
C428 a_1228_3480# VSS 0.64009f
C429 a_1012_1560# VSS 0.44974f
C430 a_796_3480# VSS 0.63814f
C431 a_580_1560# VSS 0.54364f
C432 a_364_1560# VSS 1.89817f $ **FLOATING
C433 a_3480_6364# VSS 0.59103f $ **FLOATING
C434 xa1.xa2.xa1.G VSS 15.9747f
C435 a_3480_7164# VSS 0.49536f $ **FLOATING
C436 a_3480_7432# VSS 0.05726f $ **FLOATING
C437 xa1.xa2.xd1.D VSS 3.92691f
C438 a_3480_8232# VSS 0.02588f $ **FLOATING
C439 a_15656_9218# VSS 0.48111f $ **FLOATING
C440 a_15656_9378# VSS 0.36545f $ **FLOATING
C441 xb1.xe.D VSS 1.88822f
C442 a_15656_9858# VSS 0.36516f $ **FLOATING
C443 a_15656_10018# VSS 0.48073f $ **FLOATING
C444 a_13824_9218# VSS 0.02798f $ **FLOATING
C445 xb1.xa2.P VSS 9.14989f
C446 a_13824_10018# VSS 0.09681f $ **FLOATING
C447 a_160_9538# VSS 0.02791f $ **FLOATING
C448 xa1.xb1.S VSS 10.4526f
C449 a_13824_11098# VSS 0.50256f $ **FLOATING
C450 a_13824_11258# VSS 0.4976f $ **FLOATING
C451 xb1.xb3.D VSS 12.5036f
C452 a_13824_11738# VSS 0.50771f $ **FLOATING
C453 a_13824_11898# VSS 0.5646f $ **FLOATING
C454 xa1.xe1.G VSS 19.6181f
C455 a_160_11938# VSS 0.02748f $ **FLOATING
C456 a_13824_12378# VSS 0.64355f $ **FLOATING
C457 xb3.A VSS 20.7441f
C458 a_13824_13178# VSS 0.59593f $ **FLOATING
C459 xb1.xb2.S VSS 12.8544f
.ends

