magic
tech sky130A
magscale 1 2
timestamp 1744453268
<< viali >>
rect 3289 8253 3419 8383
rect 3290 6904 3358 6972
rect 442 4273 539 4370
rect 2304 4200 2380 4440
rect 3310 2343 3409 2442
rect 3383 1481 3450 1548
rect 5223 1475 5293 1545
rect 2242 1295 2343 1396
rect -33 901 37 971
rect 3374 774 3454 854
rect 5160 -212 5388 28
<< metal1 >>
rect 3283 8389 3425 8395
rect 2622 8238 2962 8334
rect 3283 8241 3425 8247
rect 2622 8121 3024 8238
rect 3141 8121 3147 8238
rect 3608 8142 3800 8148
rect 2622 8028 2962 8121
rect 3480 8034 3544 8040
rect 3608 7994 3800 8000
rect 3480 7976 3544 7982
rect 3466 7630 3497 7722
rect 3558 7630 3564 7722
rect 3466 7574 3558 7630
rect 3992 7357 4184 7698
rect 3610 7240 3616 7357
rect 3733 7330 4184 7357
rect 4242 7330 4302 7336
rect 3733 7270 4242 7330
rect 3733 7240 4184 7270
rect 4242 7264 4302 7270
rect 3284 6978 3364 6984
rect 3284 6892 3364 6898
rect 3602 6842 3608 7034
rect 3688 6842 3694 7034
rect 3992 6954 4184 7240
rect 3480 6574 3544 6580
rect 3480 6504 3544 6510
rect 5922 4730 5928 4922
rect 6120 4730 6126 4922
rect 4693 4555 4699 4697
rect 4841 4555 4847 4697
rect 2298 4440 2386 4452
rect 436 4376 545 4382
rect 436 4261 545 4267
rect 2298 4200 2304 4440
rect 2380 4364 2386 4440
rect 2380 4322 3884 4364
rect 2380 4276 4108 4322
rect 2380 4200 2386 4276
rect 2298 4188 2386 4200
rect 3463 4141 3542 4276
rect 3785 4189 4108 4276
rect 4699 4189 4841 4555
rect 5327 4189 5409 4195
rect 3785 4148 5327 4189
rect 3457 4062 3463 4141
rect 3542 4062 3548 4141
rect 3790 4107 5327 4148
rect 3790 4036 4108 4107
rect 5327 4101 5409 4107
rect 3066 2907 3258 2908
rect 2919 2568 3655 2907
rect 2919 2520 3258 2568
rect 3304 2448 3415 2454
rect 3755 2445 3761 2539
rect 3855 2445 3861 2539
rect 3304 2331 3415 2337
rect 4096 2374 4288 2582
rect 4096 2310 4382 2374
rect 4446 2310 4452 2374
rect 3588 1910 3640 1916
rect 4096 1870 4288 2310
rect 3588 1848 3640 1854
rect 5222 1850 5228 1914
rect 5292 1858 5480 1914
rect 5292 1850 5486 1858
rect 5410 1794 5416 1850
rect 5480 1794 5486 1850
rect 5928 1824 6120 4730
rect 3377 1554 3456 1560
rect 3377 1469 3456 1475
rect 3706 1418 3712 1610
rect 3791 1418 3797 1610
rect 5217 1551 5299 1557
rect 4151 1449 4322 1531
rect 5217 1463 5299 1469
rect 5538 1414 5544 1606
rect 5626 1414 5632 1606
rect 2236 1396 2349 1408
rect 2236 1339 2242 1396
rect 339 1295 2242 1339
rect 2343 1295 2349 1396
rect 339 1248 2349 1295
rect 339 1032 430 1248
rect 2236 1166 2349 1248
rect -39 977 43 983
rect -39 889 43 895
rect 282 840 288 1032
rect 370 929 430 1032
rect 672 1138 864 1144
rect 672 1023 864 1029
rect 2236 1090 2336 1166
rect 4145 1152 4239 1155
rect 4131 1149 4239 1152
rect 4131 1125 5695 1149
rect 370 840 376 929
rect 2236 860 2349 1090
rect 4131 1065 4145 1125
rect 4239 1055 5695 1125
rect 3770 910 3846 948
rect 2236 768 2240 860
rect 2332 768 2349 860
rect 2236 574 2349 768
rect 3368 860 3460 866
rect 3368 762 3460 768
rect 3706 718 3712 910
rect 3804 776 3846 910
rect 4145 839 4239 1031
rect 5601 803 5695 1055
rect 5928 784 6120 1522
rect 3804 718 3810 776
rect 4841 742 5125 765
rect 160 356 224 486
rect 766 360 830 564
rect 2126 471 2522 574
rect 766 356 1944 360
rect 160 296 1944 356
rect 2008 296 2014 360
rect 160 292 830 296
rect 2122 276 2522 471
rect 4841 458 5482 742
rect 2578 360 2642 366
rect 2642 358 3652 360
rect 2642 298 2874 358
rect 2934 298 3652 358
rect 4841 345 5125 458
rect 4841 343 5027 345
rect 2642 296 3652 298
rect 2578 290 2642 296
rect 2168 28 2408 276
rect 5154 28 5394 40
rect 2168 -212 5160 28
rect 5388 -212 5394 28
rect 5154 -224 5394 -212
<< via1 >>
rect 3283 8383 3425 8389
rect 3283 8253 3289 8383
rect 3289 8253 3419 8383
rect 3419 8253 3425 8383
rect 3283 8247 3425 8253
rect 3024 8121 3141 8238
rect 3608 8000 3800 8142
rect 3497 7630 3558 7722
rect 3616 7240 3733 7357
rect 4242 7270 4302 7330
rect 3284 6972 3364 6978
rect 3284 6904 3290 6972
rect 3290 6904 3358 6972
rect 3358 6904 3364 6972
rect 3284 6898 3364 6904
rect 3608 6842 3688 7034
rect 3480 6510 3544 6574
rect 5928 4730 6120 4922
rect 4699 4555 4841 4697
rect 436 4370 545 4376
rect 436 4273 442 4370
rect 442 4273 539 4370
rect 539 4273 545 4370
rect 436 4267 545 4273
rect 3463 4062 3542 4141
rect 5327 4107 5409 4189
rect 3304 2442 3415 2448
rect 3761 2445 3855 2539
rect 3304 2343 3310 2442
rect 3310 2343 3409 2442
rect 3409 2343 3415 2442
rect 3304 2337 3415 2343
rect 4382 2310 4446 2374
rect 3588 1854 3640 1910
rect 5228 1850 5292 1914
rect 3377 1548 3456 1554
rect 3377 1481 3383 1548
rect 3383 1481 3450 1548
rect 3450 1481 3456 1548
rect 3377 1475 3456 1481
rect 3712 1418 3791 1610
rect 5217 1545 5299 1551
rect 5217 1475 5223 1545
rect 5223 1475 5293 1545
rect 5293 1475 5299 1545
rect 5217 1469 5299 1475
rect 5544 1414 5626 1606
rect -39 971 43 977
rect -39 901 -33 971
rect -33 901 37 971
rect 37 901 43 971
rect -39 895 43 901
rect 288 840 370 1032
rect 672 1029 864 1138
rect 4145 1031 4239 1125
rect 2240 768 2332 860
rect 3368 854 3460 860
rect 3368 774 3374 854
rect 3374 774 3454 854
rect 3454 774 3460 854
rect 3368 768 3460 774
rect 3712 718 3804 910
rect 1944 296 2008 360
rect 2578 296 2642 360
rect 2874 298 2934 358
<< metal2 >>
rect 3277 8247 3283 8389
rect 3425 8247 4841 8389
rect 3024 8238 3141 8244
rect 3633 8142 3775 8247
rect 3024 7357 3141 8121
rect 3602 8000 3608 8142
rect 3800 8000 3806 8142
rect 3497 7722 3558 7728
rect 3558 7646 3872 7707
rect 3928 7646 3937 7707
rect 3497 7624 3558 7630
rect 3616 7357 3733 7363
rect 3024 7240 3160 7357
rect 3267 7240 3616 7357
rect 4236 7270 4242 7330
rect 4302 7270 4308 7330
rect 3616 7234 3733 7240
rect 4242 7184 4302 7270
rect 4235 7128 4244 7184
rect 4300 7128 4309 7184
rect 4242 7126 4302 7128
rect 3608 7034 3688 7040
rect 3038 6898 3284 6978
rect 3364 6898 3608 6978
rect 2487 4960 2577 4962
rect 3038 4960 3118 6898
rect 3608 6836 3688 6842
rect 3474 6510 3480 6574
rect 3544 6510 3550 6574
rect 2481 4953 3119 4960
rect 2481 4863 2487 4953
rect 2577 4863 3119 4953
rect 2481 4857 3119 4863
rect 2487 4854 2577 4857
rect 430 4267 436 4376
rect 545 4267 823 4376
rect 714 1138 823 4267
rect 3038 2448 3118 4857
rect 3483 4538 3542 6510
rect 4699 4697 4841 8247
rect 5928 4922 6120 4928
rect 5919 4730 5928 4922
rect 5928 4724 6120 4730
rect 4699 4549 4841 4555
rect 3413 4462 3422 4538
rect 3478 4462 3550 4538
rect 3463 4141 3542 4147
rect 5321 4107 5327 4189
rect 5409 4107 5415 4189
rect 3038 2337 3304 2448
rect 3415 2337 3421 2448
rect 3038 2234 3152 2337
rect 288 1032 370 1038
rect -45 895 -39 977
rect 43 895 288 977
rect 666 1029 672 1138
rect 864 1029 870 1138
rect 3041 860 3152 2234
rect 3463 1554 3542 4062
rect 3761 2539 3855 2545
rect 3761 2245 3855 2445
rect 4382 2374 4446 2380
rect 3761 2151 4239 2245
rect 3588 1910 3644 1919
rect 3582 1854 3588 1910
rect 3644 1854 3646 1910
rect 3588 1845 3644 1854
rect 3712 1610 3791 1616
rect 3371 1475 3377 1554
rect 3456 1475 3712 1554
rect 3712 1412 3791 1418
rect 4145 1125 4239 2151
rect 4382 2100 4446 2310
rect 4377 2044 4386 2100
rect 4442 2044 4451 2100
rect 4382 2040 4446 2044
rect 5034 1914 5070 1926
rect 5228 1914 5292 1920
rect 5025 1850 5034 1914
rect 5090 1850 5228 1914
rect 5034 1839 5070 1850
rect 5228 1844 5292 1850
rect 5327 1551 5409 4107
rect 5544 1606 5626 1612
rect 5211 1469 5217 1551
rect 5299 1469 5544 1551
rect 5544 1408 5626 1414
rect 4139 1031 4145 1125
rect 4239 1031 4245 1125
rect 3712 910 3804 916
rect 288 834 370 840
rect 2234 768 2240 860
rect 2332 768 3368 860
rect 3460 768 3712 860
rect 3712 712 3804 718
rect 2874 586 2934 588
rect 2867 530 2876 586
rect 2932 530 2941 586
rect 1944 360 2008 366
rect 2008 296 2578 360
rect 2642 296 2648 360
rect 2874 358 2934 530
rect 1944 290 2008 296
rect 2874 292 2934 298
<< via2 >>
rect 3872 7646 3928 7707
rect 3160 7240 3267 7357
rect 4244 7128 4300 7184
rect 2487 4863 2577 4953
rect 5928 4730 6065 4922
rect 3422 4462 3478 4538
rect 3588 1854 3640 1910
rect 3640 1854 3644 1910
rect 4386 2044 4442 2100
rect 5034 1850 5090 1914
rect 2876 530 2932 586
<< metal3 >>
rect 3867 7707 3933 7712
rect 3867 7646 3872 7707
rect 3928 7646 3933 7707
rect 3867 7641 3933 7646
rect 3155 7357 3272 7362
rect 2746 7240 3160 7357
rect 3267 7240 3272 7357
rect 3155 7235 3272 7240
rect 3870 6148 3931 7641
rect 4239 7184 4305 7189
rect 4239 7128 4244 7184
rect 4300 7128 4305 7184
rect 4239 7123 4305 7128
rect 4242 7008 4302 7123
rect 4234 6944 4240 7008
rect 4304 6944 4310 7008
rect 2101 4958 2199 4963
rect 2100 4957 2582 4958
rect 2100 4859 2101 4957
rect 2199 4953 2582 4957
rect 2199 4863 2487 4953
rect 2577 4863 2582 4953
rect 2199 4859 2582 4863
rect 2100 4858 2582 4859
rect 4089 4900 4236 5513
rect 5923 4922 6070 4927
rect 5923 4900 5928 4922
rect 2101 4853 2199 4858
rect 4089 4753 5928 4900
rect 5923 4730 5928 4753
rect 6065 4730 6070 4922
rect 5923 4725 6070 4730
rect 3417 4538 3483 4543
rect 3417 4530 3422 4538
rect 2874 4470 3422 4530
rect 2874 591 2934 4470
rect 3417 4462 3422 4470
rect 3478 4462 3483 4538
rect 3417 4457 3483 4462
rect 4381 2100 4447 2105
rect 4381 2044 4386 2100
rect 4442 2044 4447 2100
rect 4381 2039 4447 2044
rect 3583 1914 3649 1915
rect 4382 1914 4446 2039
rect 5029 1914 5095 1919
rect 3583 1910 5034 1914
rect 3583 1854 3588 1910
rect 3644 1854 5034 1910
rect 3583 1850 5034 1854
rect 5090 1850 5095 1914
rect 3583 1849 3649 1850
rect 5029 1845 5095 1850
rect 2871 586 2937 591
rect 2871 530 2876 586
rect 2932 530 2937 586
rect 2871 525 2937 530
<< via3 >>
rect 4240 6944 4304 7008
rect 2101 4859 2199 4957
<< metal4 >>
rect 4239 7008 4305 7009
rect 4239 6944 4240 7008
rect 4304 6944 4305 7008
rect 4239 6943 4305 6944
rect 4242 6340 4302 6943
rect 2100 4957 2200 5420
rect 2100 4859 2101 4957
rect 2199 4859 2200 4957
rect 2100 4858 2200 4859
use JNWATR_NCH_4C5F0  xa1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 382
box -184 -128 1336 928
use JNWTR_RPPO8  xa2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1744286843
transform 1 0 0 0 1 1280
box 0 0 2744 3440
use JNWATR_NCH_4C5F0  xc1
timestamp 1740610800
transform 1 0 3424 0 1 222
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xc2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 3424 0 1 1280
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xc3
timestamp 1740610800
transform 1 0 3424 0 1 2336
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xd1
timestamp 1740610800
transform 1 0 5256 0 1 210
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xd2
timestamp 1740610800
transform 1 0 5256 0 1 1280
box -184 -128 1336 928
use JNWTR_CAPX4  xf ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1744367799
transform 1 0 -212 0 1 5320
box 480 0 3120 2640
use JNWTR_CAPX1  xg1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 3320 0 1 5320
box 0 0 1080 1080
use JNWATR_NCH_4C5F0  xg2
timestamp 1740610800
transform 1 0 3320 0 1 6386
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xg3
timestamp 1740610800
transform 1 0 3320 0 1 7454
box -184 -128 1336 928
use JNWATR_NCH_4CTAPBOT  XJNWATR_NCH_4CTAPBOT0 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 -174
box -184 -128 1336 608
use JNWATR_NCH_4CTAPBOT  XJNWATR_NCH_4CTAPBOT1
timestamp 1740610800
transform 1 0 3424 0 1 -252
box -184 -128 1336 608
use JNWATR_NCH_4CTAPBOT  XJNWATR_NCH_4CTAPBOT3
timestamp 1740610800
transform 1 0 5256 0 1 -332
box -184 -128 1336 608
use JNWATR_NCH_4CTAPTOP  XJNWATR_NCH_4CTAPTOP2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 3418 0 1 3150
box -184 -128 1336 608
use JNWATR_PCH_4CTAPTOP  XJNWATR_PCH_4CTAPTOP4 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 5256 0 1 2080
box -184 -128 1336 608
use JNWATR_PCH_4CTAPTOP  XJNWATR_PCH_4CTAPTOP5
timestamp 1740610800
transform 1 0 3320 0 1 8298
box -184 -128 1336 608
<< labels >>
flabel metal1 3798 4038 4092 4308 0 FreeSans 800 0 0 0 VDD
port 2 nsew default input
flabel metal1 2636 8044 2942 8308 0 FreeSans 800 0 0 0 Diff_Out
port 4 nsew default output
flabel metal1 2928 2532 3220 2884 0 FreeSans 800 0 0 0 V_minus
port 6 nsew default input
flabel metal1 2142 298 2516 558 0 FreeSans 800 0 0 0 VSS
port 8 nsew default input
flabel metal1 4850 350 5098 742 0 FreeSans 800 0 0 0 V_pluss
port 10 nsew default input
<< properties >>
string FIXED_BBOX 0 0 6408 8480
<< end >>
