magic
tech sky130A
magscale 1 2
timestamp 1744377898
<< viali >>
rect -39 12103 63 12205
rect -31 9321 56 9408
rect 2690 8880 2918 9120
rect 412 7712 652 7940
rect 3868 7712 4108 7940
rect 4282 6458 4510 6686
rect 410 4210 638 4438
rect 844 4200 1084 4428
rect 1326 4210 1411 4295
rect 5098 2968 5198 3068
rect 6938 1914 7031 2007
rect 5106 1435 5195 1524
rect -29 949 77 1055
rect 6924 1028 7013 1117
rect 5056 628 5248 808
<< metal1 >>
rect 2128 12250 2296 12270
rect -45 12211 69 12217
rect 131 12123 2296 12250
rect -45 12091 69 12097
rect 160 11680 228 12123
rect 306 11855 312 11880
rect 297 11741 303 11855
rect 417 11741 423 11855
rect 306 11712 312 11741
rect 426 11712 432 11880
rect 672 11090 864 11356
rect 672 11080 1628 11090
rect 672 10898 1860 11080
rect 1468 10834 1860 10898
rect 1468 10741 1695 10834
rect 1788 10741 1860 10834
rect 1468 10618 1860 10741
rect 2128 9832 2296 12123
rect 2376 10000 2568 10006
rect 2376 9802 2568 9808
rect 672 9472 864 9478
rect -37 9414 62 9420
rect -37 9309 62 9315
rect 137 8443 239 9405
rect 306 9280 312 9448
rect 411 9280 417 9448
rect 672 9373 864 9379
rect 1992 8698 2056 9348
rect 2116 9256 2122 9448
rect 2314 9256 2320 9448
rect 2684 9120 2924 9132
rect 2684 8880 2690 9120
rect 2918 9059 4802 9120
rect 2918 8945 3061 9059
rect 3175 8945 4802 9059
rect 2918 8880 4802 8945
rect 2684 8868 2924 8880
rect 1986 8634 1992 8698
rect 2056 8634 2062 8698
rect 137 8341 2039 8443
rect 400 7940 664 7946
rect 400 7712 412 7940
rect 652 7712 664 7940
rect 400 7706 664 7712
rect 412 6692 652 7706
rect 412 6452 970 6692
rect 1210 6452 1216 6692
rect 682 5988 922 5994
rect 404 5748 682 5988
rect 404 4438 644 5748
rect 682 5742 922 5748
rect 404 4210 410 4438
rect 638 4210 644 4438
rect 404 4198 644 4210
rect 832 4428 1096 4434
rect 832 4200 844 4428
rect 1084 4200 1096 4428
rect 1742 4301 1839 4307
rect 1314 4295 1742 4301
rect 1314 4210 1326 4295
rect 1411 4210 1742 4295
rect 1314 4204 1742 4210
rect 832 4194 1096 4200
rect 1742 4198 1839 4204
rect 879 1676 1050 4194
rect 683 1505 1050 1676
rect 683 1238 854 1505
rect 160 1174 854 1238
rect -35 1061 83 1067
rect -41 943 -35 1061
rect 83 943 89 1061
rect 160 1022 224 1174
rect -35 937 83 943
rect 288 918 294 1086
rect 412 918 418 1086
rect 683 923 854 1174
rect 147 153 249 449
rect 672 253 864 558
rect 1937 341 2039 8341
rect 3856 7940 4120 7946
rect 3856 7712 3868 7940
rect 4108 7712 4120 7940
rect 3856 7706 4120 7712
rect 3868 7332 4108 7706
rect 3868 7086 4108 7092
rect 2364 6692 2604 6698
rect 4562 6692 4802 8880
rect 5561 6692 6085 6791
rect 2604 6686 6085 6692
rect 2604 6458 4282 6686
rect 4510 6580 6085 6686
rect 6558 6580 6663 6586
rect 4510 6475 6558 6580
rect 4510 6458 6085 6475
rect 6558 6469 6663 6475
rect 2604 6452 6085 6458
rect 2364 6446 2604 6452
rect 4714 4301 4811 6452
rect 5490 6297 6085 6452
rect 4708 4204 4714 4301
rect 4811 4204 4817 4301
rect 5490 3102 5606 6297
rect 5092 3074 5204 3080
rect 5092 2956 5204 2962
rect 5458 2934 5464 3102
rect 5576 2960 5606 3102
rect 5824 3102 6016 3108
rect 5576 2934 5582 2960
rect 5824 2904 6016 2910
rect 5434 2678 5440 2870
rect 5558 2678 5564 2870
rect 5310 2278 5374 2462
rect 5310 2208 5374 2214
rect 4476 1978 4890 2170
rect 4476 1914 5376 1978
rect 4476 1844 4890 1914
rect 4479 1734 4890 1844
rect 5824 1828 6016 2606
rect 7144 2342 7804 2406
rect 7144 2278 7208 2342
rect 6234 2214 6240 2278
rect 6304 2214 7208 2278
rect 7740 2216 7804 2342
rect 6932 2013 7037 2019
rect 6932 1902 7037 1908
rect 7266 1864 7272 2056
rect 7377 1864 7383 2056
rect 2464 1704 3158 1706
rect 2464 1214 3268 1704
rect 5100 1530 5201 1536
rect 5100 1423 5201 1429
rect 5480 1530 5581 1536
rect 5480 1423 5581 1429
rect 2464 1121 5571 1214
rect 2464 1061 3268 1121
rect 2464 943 2587 1061
rect 2705 943 3268 1061
rect 2464 882 3268 943
rect 5056 814 5248 1121
rect 5044 808 5260 814
rect 5044 628 5056 808
rect 5248 628 5260 808
rect 5044 622 5260 628
rect 5478 624 5571 1121
rect 6918 1123 7019 1129
rect 6918 1016 7019 1022
rect 7266 976 7272 1168
rect 7373 976 7379 1168
rect 7656 1024 7848 1752
rect 5846 636 5852 737
rect 5953 636 5959 737
rect 1937 253 2043 341
rect 1941 155 2043 253
rect 1941 153 4246 155
rect 147 128 4246 153
rect 5312 128 5376 388
rect 7144 320 7208 592
rect 8374 406 8658 818
rect 8466 320 8530 406
rect 7144 256 8530 320
rect 147 64 5376 128
rect 147 53 4246 64
rect 147 51 2043 53
<< via1 >>
rect -45 12205 69 12211
rect -45 12103 -39 12205
rect -39 12103 63 12205
rect 63 12103 69 12205
rect -45 12097 69 12103
rect 303 11741 417 11855
rect 1695 10741 1788 10834
rect 2376 9808 2568 10000
rect -37 9408 62 9414
rect -37 9321 -31 9408
rect -31 9321 56 9408
rect 56 9321 62 9408
rect -37 9315 62 9321
rect 312 9280 411 9448
rect 672 9379 864 9472
rect 2122 9256 2314 9448
rect 3061 8945 3175 9059
rect 1992 8634 2056 8698
rect 970 6452 1210 6692
rect 682 5748 922 5988
rect 1742 4204 1839 4301
rect -35 1055 83 1061
rect -35 949 -29 1055
rect -29 949 77 1055
rect 77 949 83 1055
rect -35 943 83 949
rect 294 918 412 1086
rect 3868 7092 4108 7332
rect 2364 6452 2604 6692
rect 6558 6475 6663 6580
rect 4714 4204 4811 4301
rect 5092 3068 5204 3074
rect 5092 2968 5098 3068
rect 5098 2968 5198 3068
rect 5198 2968 5204 3068
rect 5092 2962 5204 2968
rect 5464 2934 5576 3102
rect 5824 2910 6016 3102
rect 5310 2214 5374 2278
rect 6240 2214 6304 2278
rect 6932 2007 7037 2013
rect 6932 1914 6938 2007
rect 6938 1914 7031 2007
rect 7031 1914 7037 2007
rect 6932 1908 7037 1914
rect 7272 1864 7377 2056
rect 5100 1524 5201 1530
rect 5100 1435 5106 1524
rect 5106 1435 5195 1524
rect 5195 1435 5201 1524
rect 5100 1429 5201 1435
rect 5480 1429 5581 1530
rect 2587 943 2705 1061
rect 6918 1117 7019 1123
rect 6918 1028 6924 1117
rect 6924 1028 7013 1117
rect 7013 1028 7019 1117
rect 6918 1022 7019 1028
rect 7272 976 7373 1168
rect 5852 636 5953 737
<< metal2 >>
rect -51 12097 -45 12211
rect 69 12097 3175 12211
rect 303 11855 417 12097
rect 303 11735 417 11741
rect 1632 10834 1715 10838
rect 1627 10829 1695 10834
rect 1627 10746 1632 10829
rect 1627 10741 1695 10746
rect 1788 10741 1794 10834
rect 1632 10737 1715 10741
rect 2376 10000 2568 10009
rect 2370 9808 2376 10000
rect 2568 9808 2574 10000
rect 672 9472 864 9481
rect 312 9448 411 9454
rect -43 9315 -37 9414
rect 62 9315 312 9414
rect 666 9379 672 9472
rect 864 9379 870 9472
rect 2122 9448 2314 9454
rect 312 8698 411 9280
rect 1992 8698 2056 8704
rect 312 8634 1992 8698
rect 312 4782 411 8634
rect 1992 8628 2056 8634
rect 2122 8522 2314 9256
rect 3061 9059 3175 12097
rect 3061 8939 3175 8945
rect 2122 8330 6016 8522
rect 3862 7092 3868 7332
rect 4108 7092 4114 7332
rect 970 6692 1210 6698
rect 1210 6452 2364 6692
rect 2604 6452 2610 6692
rect 970 6446 1210 6452
rect 3868 5988 4108 7092
rect 676 5748 682 5988
rect 922 5748 4108 5988
rect 312 4683 1575 4782
rect 294 1086 412 1092
rect -41 943 -35 1061
rect 83 943 294 1061
rect 1476 1061 1575 4683
rect 4714 4301 4811 4307
rect 1736 4204 1742 4301
rect 1839 4204 4714 4301
rect 4714 4198 4811 4204
rect 5464 3102 5576 3108
rect 5824 3102 6016 8330
rect 6552 6475 6558 6580
rect 6663 6475 6669 6580
rect 5086 2962 5092 3074
rect 5204 2962 5464 3074
rect 5464 2928 5576 2934
rect 5818 2910 5824 3102
rect 6016 2910 6022 3102
rect 6558 2833 6663 6475
rect 6561 2715 6663 2833
rect 6240 2278 6304 2284
rect 5304 2214 5310 2278
rect 5374 2214 6240 2278
rect 6240 2208 6304 2214
rect 6558 2013 6663 2715
rect 7272 2056 7377 2062
rect 6558 1908 6932 2013
rect 7037 1908 7272 2013
rect 7272 1858 7377 1864
rect 5094 1429 5100 1530
rect 5201 1429 5480 1530
rect 5581 1429 5957 1530
rect 5856 1123 5957 1429
rect 7272 1168 7373 1174
rect 412 943 2587 1061
rect 2705 943 2713 1061
rect 5852 1022 6918 1123
rect 7019 1022 7272 1123
rect 294 912 412 918
rect 5852 737 5953 1022
rect 7272 970 7373 976
rect 5852 630 5953 636
<< via2 >>
rect 1632 10746 1695 10829
rect 1695 10746 1715 10829
rect 2376 9818 2568 10000
rect 672 9389 864 9472
<< metal3 >>
rect 1556 10834 1647 10839
rect 1555 10833 1720 10834
rect 1555 10742 1556 10833
rect 1647 10829 1720 10833
rect 1715 10746 1720 10829
rect 1647 10742 1720 10746
rect 1555 10741 1720 10742
rect 1556 10736 1647 10741
rect 844 10206 2568 10398
rect 2376 10005 2568 10206
rect 2371 10000 2573 10005
rect 2371 9818 2376 10000
rect 2568 9818 2573 10000
rect 2371 9813 2573 9818
rect 667 9477 869 9483
rect 667 9380 869 9386
<< via3 >>
rect 1556 10829 1647 10833
rect 1556 10746 1632 10829
rect 1632 10746 1647 10829
rect 1556 10742 1647 10746
rect 667 9472 869 9477
rect 667 9389 672 9472
rect 672 9389 864 9472
rect 864 9389 869 9472
rect 667 9386 869 9389
<< metal4 >>
rect 722 10833 1648 10834
rect 722 10742 1556 10833
rect 1647 10742 1648 10833
rect 722 10741 1648 10742
rect 722 9478 815 10741
rect 666 9477 870 9478
rect 666 9386 667 9477
rect 869 9386 870 9477
rect 666 9385 870 9386
use JNWATR_PCH_4C1F2  xa1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 326
box -184 -128 1336 928
use JNWTR_RPPO2  xa2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1744368746
transform 1 0 0 0 1 1280
box 0 0 1448 3440
use JNWTR_RPPO16  xa3 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1744368746
transform 1 0 0 0 1 4792
box 0 0 4472 3440
use JNWATR_PCH_4C1F2  xb1
timestamp 1740610800
transform 1 0 5152 0 1 -32
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xb2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 5152 0 1 1280
box -184 -128 1336 928
use JNWATR_NCH_4C1F2  xb3 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 5152 0 1 2342
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xc2
timestamp 1740610800
transform 1 0 6984 0 1 480
box -184 -128 1336 928
use JNWATR_NCH_4C1F2  xc3
timestamp 1740610800
transform 1 0 6984 0 1 1536
box -184 -128 1336 928
use JNWATR_NCH_4C1F2  xd2
timestamp 1740610800
transform 1 0 0 0 1 11120
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  xd
timestamp 1740610800
transform 1 0 0 0 1 9240
box -184 -128 1336 928
use JNWTR_CAPX1  xd1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 0 0 1 10040
box 0 0 1080 1080
use JNWATR_NCH_2C1F2  xe ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 1832 0 1 9240
box -184 -128 1208 928
use JNWATR_NCH_2CTAPBOT  XJNWATR_NCH_2CTAPBOT7 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 1832 0 1 8760
box -184 -128 1208 608
use JNWATR_NCH_2CTAPTOP  XJNWATR_NCH_2CTAPTOP8 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 1832 0 1 10040
box -184 -128 1208 608
use JNWATR_NCH_4CTAPTOP  XJNWATR_NCH_4CTAPTOP2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 5152 0 1 3124
box -184 -128 1336 608
use JNWATR_NCH_4CTAPTOP  XJNWATR_NCH_4CTAPTOP4
timestamp 1740610800
transform 1 0 6984 0 1 2274
box -184 -128 1336 608
use JNWATR_NCH_4CTAPTOP  XJNWATR_NCH_4CTAPTOP6
timestamp 1740610800
transform 1 0 0 0 1 11920
box -184 -128 1336 608
use JNWATR_PCH_4CTAPBOT  XJNWATR_PCH_4CTAPBOT0 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 -102
box -184 -128 1336 608
use JNWATR_PCH_4CTAPBOT  XJNWATR_PCH_4CTAPBOT1
timestamp 1740610800
transform 1 0 5152 0 1 -458
box -184 -128 1336 608
use JNWATR_PCH_4CTAPBOT  XJNWATR_PCH_4CTAPBOT3
timestamp 1740610800
transform 1 0 6984 0 1 0
box -184 -128 1336 608
use JNWATR_PCH_4CTAPBOT  XJNWATR_PCH_4CTAPBOT5
timestamp 1740610800
transform 1 0 0 0 1 8760
box -184 -128 1336 608
<< labels >>
flabel metal1 5578 6322 6062 6762 0 FreeSans 800 0 0 0 VSS
port 3 nsew
flabel metal1 4488 1750 4870 2144 0 FreeSans 800 0 0 0 VIN+
port 5 nsew
flabel metal1 8388 416 8640 790 0 FreeSans 800 0 0 0 VIN-
port 7 nsew
flabel metal1 1484 10630 1850 11060 0 FreeSans 800 0 0 0 VOUT
port 9 nsew
flabel metal1 2482 894 3266 1678 0 FreeSans 800 0 0 0 VDD
port 11 nsew
<< properties >>
string FIXED_BBOX 0 0 8136 12400
<< end >>
