** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/temo_effected_current.sch
.subckt temo_effected_current VDD Vref OUT VSS
*.PININFO Vref:O VDD:I VSS:I OUT:O
xe2 Vref GATE VDD VDD JNWATR_PCH_4C5F0
xe1 LEFT_SIDE GATE VDD VDD JNWATR_PCH_4C5F0
xe3 OUT GATE VDD VDD JNWATR_PCH_4C5F0
xb1 VSS VSS LEFT_SIDE VDD JNWATR_PCH_4C5F0
xb2 VSS VSS VR VDD JNWATR_PCH_4C5F0
xc1 VR RIGHT_SIDE VSS JNWTR_RPPO2
xc2 RIGHT_SIDE Vref VSS JNWTR_RPPO8
x1 VDD LEFT_SIDE GATE RIGHT_SIDE VSS SKY_OTA
.ends

* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym # of pins=4
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sch
.subckt JNWATR_PCH_4C5F0 D G S B
*.PININFO D:B G:B S:B B:B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=3.2 nf=2 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO2.sym # of pins=3
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO2.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO2.sch
.subckt JNWTR_RPPO2 N P B
*.PININFO P:B N:B B:B
XXA1 N P B JNWTR_RES2
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO8.sym # of pins=3
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO8.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO8.sch
.subckt JNWTR_RPPO8 N P B
*.PININFO P:B N:B B:B
XXA1 N P B JNWTR_RES8
.ends


* expanding   symbol:  JNW_GR01_SKY130A/SKY_OTA.sym # of pins=5
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/SKY_OTA.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/SKY_OTA.sch
.subckt SKY_OTA VDD V_minus Diff_Out V_pluss VSS
*.PININFO VDD:I V_minus:I V_pluss:I VSS:I Diff_Out:O
xg2 Diff_Out net4 VSS VSS JNWATR_NCH_4C5F0
xc1 net3 net4 VSS VSS JNWATR_NCH_4C5F0
xa1 net4 net4 VSS VSS JNWATR_NCH_4C5F0
xc3 net1 V_minus net3 VSS JNWATR_NCH_4C5F0
xd1 net2 V_pluss net3 VSS JNWATR_NCH_4C5F0
xg3 Diff_Out net2 VDD VDD JNWATR_PCH_4C5F0
xd2 net2 net1 VDD VDD JNWATR_PCH_4C5F0
xc2 net1 net1 VDD VDD JNWATR_PCH_4C5F0
xa2 net4 VDD VSS JNWTR_RPPO8
xf Diff_Out VSS JNWTR_CAPX4
x1 net2 Diff_Out JNWTR_CAPX1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES2.sym # of pins=3
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RES2.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RES2.sch
.subckt JNWTR_RES2 N P B
*.PININFO N:B P:B B:B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 P INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES8.sym # of pins=3
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RES8.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RES8.sch
.subckt JNWTR_RES8 N P B
*.PININFO N:B P:B B:B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 INT_3 INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_4 INT_4 INT_3 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_5 INT_5 INT_4 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_6 INT_6 INT_5 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_7 P INT_6 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym # of pins=4
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sch
.subckt JNWATR_NCH_4C5F0 D G S B
*.PININFO D:B G:B S:B B:B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=3.2 nf=2 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX4.sym # of pins=2
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX4.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX4.sch
.subckt JNWTR_CAPX4 A B
*.PININFO A:B B:B
XXA1 A B JNWTR_CAPX1
XXA2 A B JNWTR_CAPX1
XXB1 A B JNWTR_CAPX1
XXB2 A B JNWTR_CAPX1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX1.sym # of pins=2
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sch
.subckt JNWTR_CAPX1 A B
*.PININFO A:B B:B
XC1 B A sky130_fd_pr__cap_mim_m3_1 W=5 L=5 m=1
.ends

.end
