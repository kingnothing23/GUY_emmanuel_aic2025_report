* NGSPICE file created from SKYOP.ext - technology: sky130A

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt SKYOP VDD VIN- VIN+ VOUT VSS
*.subckt SKYOP VSS VIN+ VIN- VOUT VDD
X0 a_796_6992# a_580_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X1 VDD xa2.P xa2.P VDD sky130_fd_pr__pfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X2 xb3.D VDD xe.D VSS sky130_fd_pr__nfet_01v8 ad=0.4704 pd=2.9 as=0.2784 ps=1.54 w=0.96 l=0.22
X3 a_3388_6992# a_3172_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X4 a_2092_6992# a_1876_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X5 a_2956_6992# a_2740_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X6 xb2.S VIN- xb3.G xb2.S sky130_fd_pr__pfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X7 xb2.S VIN+ xb3.D xb2.S sky130_fd_pr__pfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X8 a_1660_6992# a_1444_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X9 VSS xb3.G xb3.D VSS sky130_fd_pr__nfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X10 xa2.P xa2.P VDD VDD sky130_fd_pr__pfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
X11 xe.D VDD xb3.D VSS sky130_fd_pr__nfet_01v8 ad=0.2784 pd=1.54 as=0.4704 ps=2.9 w=0.96 l=0.22
X12 a_1228_6992# a_1444_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X13 xa2.P a_580_1560# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X14 VSS a_580_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X15 a_1228_6992# a_1012_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X16 VDD xa2.P VOUT VDD sky130_fd_pr__pfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X17 VDD xa2.P xb2.S VDD sky130_fd_pr__pfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X18 a_2956_6992# a_3172_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X19 VSS xb3.G xb3.G VSS sky130_fd_pr__nfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X20 a_2524_6992# a_2740_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X21 a_2524_6992# a_2308_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X22 VOUT xa2.P VDD VDD sky130_fd_pr__pfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
X23 a_2092_6992# a_2308_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X24 xa2.N a_580_1560# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X25 xb3.D xb3.G VSS VSS sky130_fd_pr__nfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
X26 xb3.G xb3.G VSS VSS sky130_fd_pr__nfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
X27 a_796_6992# a_1012_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X28 VOUT xe.D sky130_fd_pr__cap_mim_m3_1 l=5 w=5
X29 xb3.D VIN+ xb2.S xb2.S sky130_fd_pr__pfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X30 xb3.G VIN- xb2.S xb2.S sky130_fd_pr__pfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X31 xa2.N a_3604_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X32 VSS xb3.D VOUT VSS sky130_fd_pr__nfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X33 xb2.S xa2.P VDD VDD sky130_fd_pr__pfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
X34 a_3388_6992# a_3604_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X35 a_1660_6992# a_1876_5072# VSS sky130_fd_pr__res_high_po w=0.36 l=7.36
X36 VOUT xb3.D VSS VSS sky130_fd_pr__nfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
C0 a_7144_1258# a_7144_1514# 0.06279f
C1 a_160_9858# VDD 0.49339f
C2 a_160_10018# VOUT 0.01781f
C3 xb2.S a_5312_106# 0.03384f
C4 VDD VIN+ 0.07486f
C5 xb3.G a_7144_2154# 0.11839f
C6 xb3.D VOUT 0.38036f
C7 xa2.N a_3604_5072# 0.02892f
C8 VDD a_1992_9858# 0.08122f
C9 a_5312_586# xa2.P 0.08074f
C10 xa2.P a_160_9378# 0.08242f
C11 a_3172_5072# a_3604_5072# 0.14233f
C12 VIN- a_7144_458# 0.09933f
C13 VDD a_1012_5072# 0.0263f
C14 xb2.S xb3.D 0.82144f
C15 a_364_1560# VDD 0.01489f
C16 xa2.N a_1444_5072# 0.03028f
C17 a_1012_1560# a_580_1560# 0.01515f
C18 xb2.S a_5312_2058# 0.48226f
C19 xb2.S xb3.G 0.78799f
C20 xb3.G a_7144_1514# 0.03885f
C21 xb2.S a_5312_n54# 0.01206f
C22 xa2.P a_160_944# 0.11958f
C23 a_5312_3120# a_5312_2960# 0.11476f
C24 a_1228_6992# a_796_6992# 0.21349f
C25 a_160_10018# a_160_9858# 0.11476f
C26 a_160_11098# a_160_11258# 0.11476f
C27 xa2.P a_1876_5072# 0.30811f
C28 a_160_11898# xb3.D 0.0288f
C29 a_5312_586# a_5312_746# 0.11476f
C30 xa2.P a_160_464# 0.11964f
C31 VIN+ xb3.D 0.37546f
C32 a_2956_6992# a_2524_6992# 0.21349f
C33 xa2.P xe.D 0.03572f
C34 xb3.G a_7144_1674# 0.11472f
C35 a_1992_9858# xb3.D 0.05554f
C36 a_364_1560# a_580_1560# 0.01515f
C37 a_1228_6992# a_1660_6992# 0.21349f
C38 a_5312_746# a_5312_1258# 0.02844f
C39 a_5312_2058# VIN+ 0.07261f
C40 a_3388_6992# xa2.N 0.2491f
C41 a_5312_2960# a_5312_2480# 0.01174f
C42 xa2.N a_1012_5072# 0.03684f
C43 a_3388_6992# xb3.D 0.01324f
C44 a_364_1560# xa2.N 0.01537f
C45 xb3.G VIN+ 0.03975f
C46 a_1992_10018# xe.D 0.02333f
C47 a_160_9378# a_160_9218# 0.11476f
C48 xa2.P a_160_9218# 0.02164f
C49 a_7144_458# xb3.G 0.013f
C50 xb2.S a_7144_1514# 0.05316f
C51 a_7144_1674# a_7144_2154# 0.01174f
C52 a_580_5072# VDD 0.03646f
C53 a_160_464# a_160_944# 0.01174f
C54 a_160_9858# VOUT 0.03677f
C55 a_160_11258# xb3.D 0.08168f
C56 a_160_11898# VOUT 0.01258f
C57 xa2.N a_4036_5072# 0.1466f
C58 a_5312_586# VDD 0.49275f
C59 a_160_9378# VDD 0.50229f
C60 xa2.P VDD 8.41183f
C61 xa2.P a_160_1104# 0.07112f
C62 a_160_11738# xb3.D 0.08445f
C63 a_5312_1258# VDD 0.02387f
C64 a_2956_6992# xb3.D 0.01324f
C65 xb2.S VIN+ 2.58213f
C66 a_7144_1674# a_7144_1514# 0.11476f
C67 a_5312_3120# xb3.D 0.02778f
C68 xa2.P a_2308_5072# 0.01443f
C69 xa2.P a_2092_6992# 0.12598f
C70 a_7144_458# xb2.S 0.6232f
C71 xa2.P a_160_304# 0.05442f
C72 a_1012_5072# a_1444_5072# 0.14233f
C73 VDD a_160_944# 0.50687f
C74 a_160_1104# a_160_944# 0.11476f
C75 a_160_11258# VOUT 0.03724f
C76 a_5312_2320# xb3.D 0.03393f
C77 a_4036_5072# a_3604_5072# 0.01515f
C78 a_5312_586# a_5312_106# 0.01174f
C79 a_580_5072# xa2.N 0.21356f
C80 a_364_1560# a_1012_1560# 0.06667f
C81 xa2.P a_5312_106# 0.08182f
C82 xa2.P a_580_1560# 0.22449f
C83 a_5312_2480# xb3.D 0.03329f
C84 a_5312_746# VDD 0.42427f
C85 a_5312_2320# a_5312_2058# 0.06106f
C86 VDD a_160_464# 0.50483f
C87 a_160_11738# VOUT 0.03418f
C88 a_5312_2320# xb3.G 0.02601f
C89 VDD xe.D 0.44881f
C90 xa2.P xa2.N 0.58692f
C91 xa2.P xb3.D 0.03016f
C92 a_1992_9378# xe.D 0.02838f
C93 xb3.G a_5312_2480# 0.08513f
C94 a_2308_5072# a_1876_5072# 0.14233f
C95 a_160_11098# xe.D 0.03109f
C96 a_5312_1258# xb3.D 0.013f
C97 a_580_5072# a_364_5072# 0.01515f
C98 VDD a_160_9218# 0.56296f
C99 a_1992_10018# xb3.D 0.0371f
C100 a_160_464# a_160_304# 0.11476f
C101 xe.D a_1992_9218# 0.01169f
C102 a_7144_2314# xb3.G 0.05596f
C103 VDD a_160_1104# 0.41416f
C104 VIN- VDD 0.02736f
C105 xb2.S a_5312_2320# 0.04804f
C106 a_160_11738# a_160_11898# 0.11476f
C107 a_1992_9378# VDD 0.08135f
C108 a_1876_5072# xa2.N 0.0171f
C109 a_7144_2314# a_7144_2154# 0.11476f
C110 a_160_9378# VOUT 0.03203f
C111 xa2.P VOUT 0.21783f
C112 xa2.P a_1660_6992# 0.23404f
C113 a_160_10018# xe.D 0.03583f
C114 a_5312_586# xb2.S 0.03571f
C115 xe.D xb3.D 0.79739f
C116 VDD a_1992_9218# 0.01578f
C117 xa2.P xb2.S 0.18817f
C118 VIN- a_7144_1258# 0.071f
C119 xa2.P a_1228_6992# 0.01614f
C120 VDD a_160_304# 0.58222f
C121 xa2.P a_1444_5072# 0.02072f
C122 a_1992_9378# a_1992_9218# 0.0971f
C123 a_2092_6992# a_2524_6992# 0.21349f
C124 xb2.S a_5312_1258# 0.50479f
C125 a_3388_6992# a_2956_6992# 0.21349f
C126 xa2.P a_1012_1560# 0.245f
C127 a_5312_2960# xb3.D 0.02933f
C128 a_5312_106# VDD 0.50265f
C129 VDD a_580_1560# 0.01455f
C130 a_2308_5072# a_2740_5072# 0.14233f
C131 a_160_11738# a_160_11258# 0.01174f
C132 xb3.G a_5312_2960# 0.08185f
C133 a_160_10018# VDD 0.40658f
C134 a_160_9858# a_160_9378# 0.01174f
C135 xa2.P a_160_9858# 0.08107f
C136 VDD xa2.N 0.87608f
C137 VDD xb3.D 0.56034f
C138 a_1992_9378# xb3.D 0.05643f
C139 a_1876_5072# a_1444_5072# 0.14233f
C140 a_160_10018# a_160_11098# 0.01285f
C141 xe.D VOUT 2.99968f
C142 xb3.D a_2524_6992# 0.01324f
C143 a_580_5072# a_1012_5072# 0.14233f
C144 xb2.S a_5312_746# 0.03533f
C145 VIN- xb3.G 0.44181f
C146 a_2308_5072# xa2.N 0.02767f
C147 a_2092_6992# xb3.D 0.01142f
C148 a_5312_1258# VIN+ 0.07043f
C149 xb3.D a_1992_9218# 0.02923f
C150 VOUT a_160_9218# 0.01478f
C151 xa2.P a_364_1560# 0.04127f
C152 a_364_5072# VDD 0.08277f
C153 VDD a_5312_n54# 0.58137f
C154 a_1992_10018# a_1992_9858# 0.0971f
C155 xa2.N a_2740_5072# 0.02767f
C156 VDD a_796_6992# 0.0269f
C157 a_3172_5072# a_2740_5072# 0.14233f
C158 xb3.G a_7144_1258# 0.03814f
C159 VDD VOUT 0.99117f
C160 xb2.S VDD 1.16666f
C161 VDD a_1228_6992# 0.01333f
C162 a_160_11098# VOUT 0.04366f
C163 VIN- xb2.S 3.25396f
C164 xa2.N xb3.D 0.02365f
C165 VDD a_1444_5072# 0.01168f
C166 xa2.N a_3172_5072# 0.02767f
C167 a_5312_2058# xb3.D 0.03695f
C168 xe.D a_1992_9858# 0.02992f
C169 VDD a_1012_1560# 0.02973f
C170 a_2092_6992# a_1660_6992# 0.21349f
C171 xb3.G xb3.D 0.43731f
C172 a_5312_106# a_5312_n54# 0.11476f
C173 xb2.S a_7144_1258# 0.4835f
C174 a_5312_2058# xb3.G 0.01323f
C175 a_5312_2320# a_5312_2480# 0.11476f
C176 a_364_5072# xa2.N 0.10537f
C177 VIN- VSS 0.80129f
C178 VIN+ VSS 0.71565f
C179 VOUT VSS 2.75355f
C180 VDD VSS 30.3698f
C181 a_7144_458# VSS 0.02653f $ **FLOATING
C182 a_5312_n54# VSS 0.02916f $ **FLOATING
C183 a_5312_746# VSS 0.07212f $ **FLOATING
C184 a_160_304# VSS 0.02981f $ **FLOATING
C185 a_7144_1258# VSS 0.05294f $ **FLOATING
C186 a_160_1104# VSS 0.13937f $ **FLOATING
C187 a_5312_1258# VSS 0.07213f $ **FLOATING
C188 a_7144_1514# VSS 0.41005f $ **FLOATING
C189 a_7144_1674# VSS 0.49626f $ **FLOATING
C190 a_5312_2058# VSS 0.05665f $ **FLOATING
C191 a_7144_2154# VSS 0.50871f $ **FLOATING
C192 a_7144_2314# VSS 0.61822f $ **FLOATING
C193 a_5312_2320# VSS 0.41618f $ **FLOATING
C194 a_5312_2480# VSS 0.49887f $ **FLOATING
C195 xb3.G VSS 5.61207f
C196 a_5312_2960# VSS 0.50822f $ **FLOATING
C197 a_5312_3120# VSS 0.60866f $ **FLOATING
C198 a_1012_1560# VSS 1.82365f $ **FLOATING
C199 a_580_1560# VSS 0.62373f
C200 a_364_1560# VSS 1.82183f $ **FLOATING
C201 a_4036_5072# VSS 1.99287f $ **FLOATING
C202 xa2.N VSS 5.04286f
C203 a_3604_5072# VSS 0.5397f
C204 a_3388_6992# VSS 0.64011f
C205 a_3172_5072# VSS 0.44449f
C206 a_2956_6992# VSS 0.63998f
C207 a_2740_5072# VSS 0.44331f
C208 a_2524_6992# VSS 0.63914f
C209 a_2308_5072# VSS 0.44299f
C210 a_2092_6992# VSS 0.6436f
C211 a_1876_5072# VSS 0.43952f
C212 a_1660_6992# VSS 0.64541f
C213 a_1444_5072# VSS 0.43888f
C214 a_1228_6992# VSS 0.64995f
C215 a_1012_5072# VSS 0.43635f
C216 a_796_6992# VSS 0.89975f
C217 a_580_5072# VSS 0.53141f
C218 a_364_5072# VSS 2.01377f $ **FLOATING
C219 a_1992_9218# VSS 0.48111f $ **FLOATING
C220 a_1992_9378# VSS 0.36545f $ **FLOATING
C221 xe.D VSS 2.19519f
C222 a_1992_9858# VSS 0.36516f $ **FLOATING
C223 a_1992_10018# VSS 0.48073f $ **FLOATING
C224 a_160_9218# VSS 0.02798f $ **FLOATING
C225 xa2.P VSS 9.1557f
C226 a_160_10018# VSS 0.09702f $ **FLOATING
C227 a_160_11098# VSS 0.50235f $ **FLOATING
C228 a_160_11258# VSS 0.4976f $ **FLOATING
C229 xb3.D VSS 12.5979f
C230 a_160_11738# VSS 0.50705f $ **FLOATING
C231 a_160_11898# VSS 0.5938f $ **FLOATING
C232 xb2.S VSS 12.8545f
.ends

