magic
tech sky130A
magscale 1 2
timestamp 1744453268
<< locali >>
rect 9153 120 9562 126
rect 9153 15 9159 120
rect 9264 15 9562 120
rect 9153 9 9562 15
<< viali >>
rect 294 9198 474 9378
rect 9324 6458 9552 6686
rect 12744 6468 12984 6696
rect 10523 3553 10628 3658
rect 9338 2978 9518 3158
rect 9750 2932 9990 3160
rect 7006 2200 7234 2440
rect 9159 15 9264 120
<< metal1 >>
rect 2642 11520 3238 11528
rect 2642 11486 3604 11520
rect 160 10244 224 11264
rect 288 10056 480 11482
rect 672 11294 3604 11486
rect 2642 10920 3604 11294
rect 672 10626 1670 10866
rect 160 8248 224 9700
rect 288 9378 480 9864
rect 288 9198 294 9378
rect 474 9198 480 9378
rect 669 9307 824 9783
rect 1430 9628 1670 10626
rect 2666 9838 3644 10440
rect 2666 9828 2858 9838
rect 3014 9628 3254 9838
rect 1430 9388 5162 9628
rect 288 8964 480 9198
rect 663 9152 669 9307
rect 824 9152 830 9307
rect 288 8766 480 8772
rect 160 8184 2774 8248
rect 4922 7306 5162 9388
rect 4922 7066 12984 7306
rect 12744 6702 12984 7066
rect 9318 6686 9558 6698
rect 9318 6458 9324 6686
rect 9552 6458 9558 6686
rect 12732 6696 12996 6702
rect 12732 6468 12744 6696
rect 12984 6468 12996 6696
rect 12732 6462 12996 6468
rect 9318 5384 9558 6458
rect 7376 5099 8342 5202
rect 9318 5144 9990 5384
rect 7376 4957 7449 5099
rect 7591 4957 8342 5099
rect 7376 4916 8342 4957
rect 7000 4676 8342 4916
rect 4653 4000 4808 4006
rect 3035 3845 4653 4000
rect 3035 2687 3190 3845
rect 4653 3839 4808 3845
rect 7000 2440 7240 4676
rect 7376 4668 8342 4676
rect 9750 3636 9990 5144
rect 10517 3658 10634 3670
rect 9744 3396 9750 3636
rect 9990 3396 9996 3636
rect 10517 3553 10523 3658
rect 10628 3553 10634 3658
rect 9750 3166 9990 3396
rect 7000 2200 7006 2440
rect 7234 2200 7240 2440
rect 7000 2188 7240 2200
rect 7376 3158 9530 3164
rect 7376 2978 9338 3158
rect 9518 2978 9530 3158
rect 7376 2972 9530 2978
rect 9738 3160 10002 3166
rect 7376 1706 7568 2972
rect 9738 2932 9750 3160
rect 9990 2932 10002 3160
rect 9738 2926 10002 2932
rect 7248 1150 7312 1392
rect 7760 1044 7952 1524
rect 4852 514 4858 702
rect 5046 514 5052 702
rect 7370 628 7376 820
rect 7531 628 7537 820
rect 4914 22 7102 28
rect 7248 22 7312 604
rect 7760 22 7952 712
rect 9153 120 9270 132
rect 4914 -100 8328 22
rect 9153 15 9159 120
rect 9264 15 9270 120
rect 9153 -100 9270 15
rect 10517 -100 10634 3553
rect 4914 -212 10634 -100
rect 6946 -217 10634 -212
rect 6946 -340 8332 -217
<< via1 >>
rect 669 9152 824 9307
rect 288 8772 480 8964
rect 7449 4957 7591 5099
rect 4653 3845 4808 4000
rect 9750 3396 9990 3636
rect 4858 514 5046 702
rect 7376 628 7531 820
<< metal2 >>
rect 669 9307 824 9313
rect 669 9146 824 9152
rect 282 8772 288 8964
rect 480 8772 4834 8964
rect 4642 8200 4834 8772
rect 4699 4957 7449 5099
rect 7591 4957 7597 5099
rect 4940 4000 5085 4004
rect 4647 3845 4653 4000
rect 4808 3995 5090 4000
rect 4808 3850 4940 3995
rect 5085 3850 5090 3995
rect 4808 3845 5090 3850
rect 4940 3841 5085 3845
rect 9750 3636 9990 3642
rect 9199 3396 9208 3636
rect 9438 3396 9750 3636
rect 9750 3390 9990 3396
rect 4858 3259 5046 3264
rect 4854 3081 4863 3259
rect 5041 3081 5050 3259
rect 4858 702 5046 3081
rect 7376 820 7531 826
rect 7367 628 7376 820
rect 7376 622 7531 628
rect 4858 508 5046 514
<< via2 >>
rect 674 9157 819 9302
rect 4940 3850 5085 3995
rect 9208 3396 9438 3636
rect 4863 3081 5041 3259
rect 7376 628 7521 820
<< metal3 >>
rect 669 9302 6846 9307
rect 669 9157 674 9302
rect 819 9157 6846 9302
rect 669 9152 6846 9157
rect 6691 4000 6846 9152
rect 4935 3995 6846 4000
rect 4935 3850 4940 3995
rect 5085 3850 6846 3995
rect 4935 3845 6846 3850
rect 4828 3398 4834 3635
rect 5071 3398 5077 3635
rect 4858 3259 5046 3398
rect 4858 3081 4863 3259
rect 5041 3081 5046 3259
rect 4858 3076 5046 3081
rect 6691 802 6846 3845
rect 9203 3636 9443 3641
rect 8442 3396 8448 3636
rect 8686 3396 9208 3636
rect 9438 3396 9443 3636
rect 9203 3391 9443 3396
rect 7371 820 7526 825
rect 7371 802 7376 820
rect 6691 647 7376 802
rect 7371 628 7376 647
rect 7521 628 7526 820
rect 7371 623 7526 628
<< via3 >>
rect 4834 3398 5071 3635
rect 8448 3396 8686 3636
<< metal4 >>
rect 8447 3636 8687 3637
rect 4833 3635 8448 3636
rect 4833 3398 4834 3635
rect 5071 3398 8448 3635
rect 4833 3397 8448 3398
rect 8447 3396 8448 3397
rect 8686 3396 8687 3636
rect 8447 3395 8687 3396
use SKY_OTA  xa3 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_GR01_SKY130A
timestamp 1744453268
transform 1 0 0 0 1 0
box -184 -460 6592 8906
use JNWATR_PCH_4C5F0  xb1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 7088 0 1 480
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xb2
timestamp 1740610800
transform 1 0 7088 0 1 1280
box -184 -128 1336 928
use JNWTR_RPPO2  xc1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1744368746
transform 1 0 8920 0 1 0
box 0 0 1448 3440
use JNWTR_RPPO16  xc2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1744368746
transform 1 0 8920 0 1 3536
box 0 0 4472 3440
use JNWATR_PCH_4C5F0  xe1
timestamp 1740610800
transform 1 0 0 0 1 9560
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xe2
timestamp 1740610800
transform 1 0 0 0 1 10360
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  xe3
timestamp 1740610800
transform 1 0 0 0 1 11160
box -184 -128 1336 928
use JNWATR_PCH_4CTAPBOT  XJNWATR_PCH_4CTAPBOT0 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 7088 0 1 0
box -184 -128 1336 608
use JNWATR_PCH_4CTAPBOT  XJNWATR_PCH_4CTAPBOT2
timestamp 1740610800
transform 1 0 0 0 1 9080
box -184 -128 1336 608
use JNWATR_PCH_4CTAPTOP  XJNWATR_PCH_4CTAPTOP1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 7088 0 1 2080
box -184 -128 1336 608
use JNWATR_PCH_4CTAPTOP  XJNWATR_PCH_4CTAPTOP3
timestamp 1740610800
transform 1 0 0 0 1 11960
box -184 -128 1336 608
<< labels >>
flabel metal1 6972 -304 8296 -14 0 FreeSans 800 0 0 0 VSS
port 1 nsew
flabel metal1 7416 4702 8304 5164 0 FreeSans 800 0 0 0 VDD
port 3 nsew
flabel metal1 2692 10954 3576 11496 0 FreeSans 800 0 0 0 OUT
port 5 nsew
flabel metal1 2682 9844 3624 10410 0 FreeSans 800 0 0 0 Vref
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 13392 12440
<< end >>
