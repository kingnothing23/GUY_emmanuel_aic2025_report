* NGSPICE file created from JNW_GR01.ext - technology: sky130A

.subckt JNWTR_CAPX1 A B
X0 B A sky130_fd_pr__cap_mim_m3_1 l=5 w=5
.ends

.subckt JNWATR_NCH_4C1F2 D G S B a_1056_n40#
X0 S G D B sky130_fd_pr__nfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X1 D G S B sky130_fd_pr__nfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
.ends

.subckt JNWATR_PCH_4C5F0 D G S B a_160_778# a_160_n22#
X0 S G D B sky130_fd_pr__pfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
X1 D G S B sky130_fd_pr__pfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
.ends

.subckt JNWATR_PCH_4C1F2 D G S B
X0 S G D B sky130_fd_pr__pfet_01v8 ad=0.784 pd=4.18 as=0.464 ps=2.18 w=1.6 l=0.22
X1 D G S B sky130_fd_pr__pfet_01v8 ad=0.464 pd=2.18 as=0.784 ps=4.18 w=1.6 l=0.22
.ends

.subckt JNWTR_RES2 N P 0
X0 N a_180_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X1 P a_180_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
.ends

.subckt JNWTR_RPPO2 P N B
XXA1 N P B JNWTR_RES2
.ends

.subckt JNWTR_RES16 N P 0
X0 a_2556_1800# a_2340_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X1 a_1260_1800# a_1476_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X2 a_396_1800# a_612_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X3 a_2556_1800# a_2772_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X4 a_1692_1800# a_1476_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X5 a_828_1800# a_612_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X6 a_2988_1800# a_2772_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X7 N a_180_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X8 a_2988_1800# a_3204_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X9 a_2124_1800# a_1908_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X10 a_828_1800# a_1044_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X11 a_1692_1800# a_1908_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X12 a_396_1800# a_180_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X13 P a_3204_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X14 a_2124_1800# a_2340_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X15 a_1260_1800# a_1044_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
.ends

.subckt JNWTR_RPPO16 P N B
XXA1 N P B JNWTR_RES16
.ends

.subckt JNWATR_NCH_2C1F2 D G S B a_928_n40#
X0 S G D B sky130_fd_pr__nfet_01v8 ad=0.4704 pd=2.9 as=0.2784 ps=1.54 w=0.96 l=0.22
X1 D G S B sky130_fd_pr__nfet_01v8 ad=0.2784 pd=1.54 as=0.4704 ps=2.9 w=0.96 l=0.22
.ends

.subckt SKYOP VSS VIN+ VIN- VOUT VDD
Xxd1 xe/D VOUT JNWTR_CAPX1
Xxd2 VOUT xe/S VSS VSS VSS JNWATR_NCH_4C1F2
Xxc2 xc3/G VIN- xc2/S xc2/S xc2/a_160_778# xc2/a_160_n22# JNWATR_PCH_4C5F0
Xxb1 xc2/S xd/G VDD VDD JNWATR_PCH_4C1F2
Xxc3 xc3/G xc3/G VSS VSS xc3/a_1056_n40# JNWATR_NCH_4C1F2
Xxb2 xe/S VIN+ xc2/S xc2/S xb2/a_160_778# xb2/a_160_n22# JNWATR_PCH_4C5F0
Xxa1 xd/G xd/G VDD VDD JNWATR_PCH_4C1F2
Xxb3 xe/S xc3/G VSS VSS VSS JNWATR_NCH_4C1F2
Xxa2 xd/G xa3/P VSS JNWTR_RPPO2
Xxa3 xa3/P VSS VSS JNWTR_RPPO16
Xxd VOUT xd/G VDD VDD JNWATR_PCH_4C1F2
Xxe xe/D VDD xe/S VSS VSS JNWATR_NCH_2C1F2
.ends

.subckt JNWTR_RES8 N P 0
X0 a_1260_1800# a_1476_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X1 a_396_1800# a_612_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X2 P a_1476_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X3 a_828_1800# a_612_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X4 N a_180_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X5 a_828_1800# a_1044_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X6 a_396_1800# a_180_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
X7 a_1260_1800# a_1044_n120# 0 sky130_fd_pr__res_high_po w=0.36 l=7.36
.ends

.subckt JNWTR_RPPO8 P N B
XXA1 N P B JNWTR_RES8
.ends

.subckt JNWATR_NCH_4C5F0 D G S B a_1056_n40#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.528 pd=2.26 as=0.848 ps=4.26 w=1.6 l=0.94
X1 S G D B sky130_fd_pr__nfet_01v8 ad=0.848 pd=4.26 as=0.528 ps=2.26 w=1.6 l=0.94
.ends

.subckt JNWTR_CAPX4 A B
XXB1 A B JNWTR_CAPX1
XXA1 A B JNWTR_CAPX1
XXB2 A B JNWTR_CAPX1
XXA2 A B JNWTR_CAPX1
.ends

.subckt SKY_OTA VDD Diff_Out V_minus V_pluss VSS
Xxg1 xg3/G Diff_Out JNWTR_CAPX1
Xxg2 Diff_Out xg2/G VSS VSS xg2/a_1056_n40# JNWATR_NCH_4C5F0
Xxg3 Diff_Out xg3/G VDD VDD xg3/a_160_778# xg3/a_160_n22# JNWATR_PCH_4C5F0
Xxd1 xg3/G V_pluss xd1/S VSS VSS JNWATR_NCH_4C5F0
Xxd2 xg3/G xd2/G VDD VDD xd2/a_160_778# xd2/a_160_n22# JNWATR_PCH_4C5F0
Xxc2 xd2/G xd2/G VDD VDD xc2/a_160_778# xc2/a_160_n22# JNWATR_PCH_4C5F0
Xxc1 xd1/S xg2/G VSS VSS VSS JNWATR_NCH_4C5F0
Xxc3 xd2/G V_minus xd1/S VSS VSS JNWATR_NCH_4C5F0
Xxa1 xg2/G xg2/G VSS VSS VSS JNWATR_NCH_4C5F0
Xxa2 VDD xg2/G VSS JNWTR_RPPO8
Xxf Diff_Out VSS JNWTR_CAPX4
.ends

.subckt temo_effected_current VDD VSS Vref OUT
Xxe1 xe1/D xe3/G VDD VDD xe2/a_160_n22# xe1/a_160_n22# JNWATR_PCH_4C5F0
Xxe2 Vref xe3/G VDD VDD xe3/a_160_n22# xe2/a_160_n22# JNWATR_PCH_4C5F0
Xxe3 OUT xe3/G VDD VDD xe3/a_160_778# xe3/a_160_n22# JNWATR_PCH_4C5F0
Xxc2 Vref xc2/N VSS JNWTR_RPPO8
Xxc1 xc2/N xc1/N VSS JNWTR_RPPO2
Xxb1 VSS VSS xe1/D VDD xb2/a_160_n22# xb1/a_160_n22# JNWATR_PCH_4C5F0
Xxb2 VSS VSS xc1/N VDD xb2/a_160_778# xb2/a_160_n22# JNWATR_PCH_4C5F0
Xxa2 VDD xe3/G xe1/D xc2/N VSS SKY_OTA
.ends

.subckt JNW_GR01 VDD VSS reset cmp vref
Xxb1 VSS xb3/A vref cmp VDD SKYOP
Xxa1 VDD VSS vref xb3/A temo_effected_current
Xxb2 xb3/A reset VSS VSS xb2/a_1056_n40# JNWATR_NCH_4C5F0
Xxb3 xb3/A VSS JNWTR_CAPX1
.ends

