magic
tech sky130A
magscale 1 2
timestamp 1744459438
<< viali >>
rect 13631 12527 13725 12621
<< metal1 >>
rect 5406 13749 6914 13894
rect 4089 12959 6914 13749
rect 2473 11378 2479 11950
rect 2828 11378 2834 11950
rect 4089 10992 4879 12959
rect 5406 12490 6914 12959
rect 7878 12533 9884 13802
rect 10806 12996 12002 13438
rect 10806 12932 13888 12996
rect 10806 12580 12002 12932
rect 14336 12768 14528 12774
rect 7854 12312 9884 12533
rect 10792 12412 12002 12580
rect 13625 12627 13731 12633
rect 13625 12515 13731 12521
rect 13952 12618 14144 12624
rect 14336 12618 14528 12624
rect 13952 12506 14144 12512
rect 8955 11080 9201 12312
rect 4089 10779 6388 10992
rect 8955 10834 15419 11080
rect 4089 10490 4879 10779
rect 6175 8771 6388 10779
rect 6169 8558 6175 8771
rect 6388 8558 6394 8771
rect 7305 6438 7311 6962
rect 7584 6438 7590 6962
rect 12425 6548 12431 6575
rect 12046 6302 12431 6548
rect 12704 6548 12710 6575
rect 12704 6302 13144 6548
rect 12046 5492 13144 6302
rect 12112 5482 13144 5492
rect 12869 5127 13072 5482
rect 12018 4742 12024 4982
rect 12264 4742 12270 4982
rect 12863 4924 12869 5127
rect 13072 4924 13078 5127
rect 12024 4592 12264 4742
rect 11936 4450 13328 4592
rect 11936 3318 13340 4450
rect 11980 -121 12131 3318
rect 18203 2801 18209 3039
rect 18447 2801 18453 3039
rect 18209 1899 18447 2801
rect 22055 1846 22061 2059
rect 22274 1846 22280 2059
rect 16128 1706 16773 1712
rect 16128 1497 16773 1503
rect 22061 536 22274 1846
rect 9172 -272 12131 -121
<< via1 >>
rect 2479 11378 2828 11950
rect 13625 12621 13731 12627
rect 14336 12624 14528 12768
rect 13625 12527 13631 12621
rect 13631 12527 13725 12621
rect 13725 12527 13731 12621
rect 13625 12521 13731 12527
rect 13952 12512 14144 12618
rect 6175 8558 6388 8771
rect 7311 6438 7584 6962
rect 12431 6302 12704 6575
rect 12024 4742 12264 4982
rect 12869 4924 13072 5127
rect 18209 2801 18447 3039
rect 22061 1846 22274 2059
rect 16128 1503 16773 1706
<< metal2 >>
rect 14336 12768 14528 12777
rect 13619 12521 13625 12627
rect 13731 12618 14101 12627
rect 14330 12624 14336 12768
rect 14528 12624 14534 12768
rect 13731 12521 13952 12618
rect 13946 12512 13952 12521
rect 14144 12512 14150 12618
rect 13995 12103 14101 12512
rect 2479 11950 2828 11956
rect 2828 11378 2837 11950
rect 2479 11372 2828 11378
rect 6175 8771 6388 8777
rect 6388 8558 6397 8771
rect 6175 8552 6388 8558
rect 7311 6962 7584 6968
rect 7584 6575 12704 6837
rect 7584 6564 12431 6575
rect 7311 6432 7584 6438
rect 15211 6452 15220 6692
rect 15450 6452 15459 6692
rect 12431 6296 12704 6302
rect 12024 5249 12264 5254
rect 12020 5019 12029 5249
rect 12259 5019 12268 5249
rect 12869 5127 13072 5133
rect 12024 4982 12264 5019
rect 12865 4924 12869 4936
rect 13072 4924 13076 4936
rect 12865 4743 12874 4924
rect 13067 4743 13076 4924
rect 12024 4736 12264 4742
rect 12869 4738 13072 4743
rect 18209 4028 18447 4033
rect 18205 3800 18214 4028
rect 18442 3800 18451 4028
rect 18209 3039 18447 3800
rect 22061 3162 22274 3167
rect 22057 2959 22066 3162
rect 22269 2959 22278 3162
rect 18209 2795 18447 2801
rect 22061 2059 22274 2959
rect 22061 1840 22274 1846
rect 16128 1706 16773 1715
rect 16122 1503 16128 1706
rect 16773 1503 16779 1706
<< via2 >>
rect 14336 12634 14528 12768
rect 13995 12521 14101 12617
rect 2489 11378 2828 11950
rect 6185 8558 6388 8771
rect 15220 6452 15450 6692
rect 12029 5019 12259 5249
rect 12874 4924 13067 4936
rect 12874 4743 13067 4924
rect 18214 3800 18442 4028
rect 22066 2959 22269 3162
rect 16128 1513 16773 1706
<< metal3 >>
rect 12599 13746 14068 13802
rect 18209 13746 18447 13750
rect 12599 13744 18447 13746
rect 12599 13508 18209 13744
rect 12599 13453 14068 13508
rect 18209 13502 18447 13508
rect 2484 11950 2833 11955
rect 2484 11378 2489 11950
rect 2828 11839 2833 11950
rect 12599 11839 12948 13453
rect 14360 12773 14504 13448
rect 14331 12768 14533 12773
rect 14331 12634 14336 12768
rect 14528 12634 14533 12768
rect 14331 12629 14533 12634
rect 13990 12622 14106 12628
rect 13990 12512 14106 12518
rect 2828 11490 12948 11839
rect 2828 11378 2833 11490
rect 2484 11373 2833 11378
rect 6180 8771 6393 8776
rect 6180 8558 6185 8771
rect 6388 8558 21166 8771
rect 6180 8553 6393 8558
rect 18209 8078 18447 8079
rect 18204 7842 18210 8078
rect 18446 7842 18452 8078
rect 15215 6692 15455 6697
rect 12024 6452 15220 6692
rect 15450 6452 15455 6692
rect 12024 5249 12264 6452
rect 15215 6447 15455 6452
rect 12024 5019 12029 5249
rect 12259 5019 12264 5249
rect 12024 5014 12264 5019
rect 12869 4936 13072 4941
rect 12869 4743 12874 4936
rect 13067 4743 13072 4936
rect 12869 1997 13072 4743
rect 18209 4028 18447 7842
rect 18209 3800 18214 4028
rect 18442 3800 18447 4028
rect 18209 3795 18447 3800
rect 20953 3167 21166 8558
rect 20953 3162 22274 3167
rect 20953 2959 22066 3162
rect 22269 2959 22274 3162
rect 20953 2954 22274 2959
rect 12869 1794 16552 1997
rect 16349 1711 16552 1794
rect 16123 1706 16778 1711
rect 16123 1513 16128 1706
rect 16773 1513 16778 1706
rect 16123 1508 16778 1513
<< via3 >>
rect 18209 13508 18447 13744
rect 13990 12617 14106 12622
rect 13990 12521 13995 12617
rect 13995 12521 14101 12617
rect 14101 12521 14106 12617
rect 13990 12518 14106 12521
rect 18210 7842 18446 8078
<< metal4 >>
rect 18208 13744 18448 13745
rect 18208 13508 18209 13744
rect 18447 13508 18448 13744
rect 18208 13507 18448 13508
rect 13995 12623 14101 13485
rect 13989 12622 14107 12623
rect 13989 12518 13990 12622
rect 14106 12518 14107 12622
rect 13989 12517 14107 12518
rect 18209 8078 18447 13507
rect 18209 7842 18210 8078
rect 18446 7842 18447 8078
rect 18209 7841 18447 7842
use temo_effected_current  xa1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_GR01_SKY130A
timestamp 1744454117
transform 1 0 0 0 1 0
box -184 -460 11664 12568
use SKYOP  xb1 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_GR01_SKY130A
timestamp 1744377898
transform 1 0 13664 0 1 0
box -184 -586 8658 12528
use JNWATR_NCH_4C5F0  xb2 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 13664 0 1 12400
box -184 -128 1336 928
use JNWTR_CAPX1  xb3 ~/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 13664 0 1 13200
box 0 0 1080 1080
<< labels >>
flabel metal1 12100 5494 13100 6536 0 FreeSans 1600 0 0 0 VDD
port 1 nsew default input
flabel metal1 12002 3374 13176 4504 0 FreeSans 1600 0 0 0 VSS
port 2 nsew default input
flabel metal1 10810 12452 11970 13372 0 FreeSans 1600 0 0 0 reset
port 3 nsew default input
flabel metal1 7952 12380 9844 13726 0 FreeSans 1600 0 0 0 cmp
port 4 nsew default output
flabel metal1 5458 12566 6850 13854 0 FreeSans 1600 0 0 0 vref
port 5 nsew default output
<< properties >>
string FIXED_BBOX 0 0 21800 14280
<< end >>
