** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_GR01_SKY130A/SKYOP.sch
.subckt SKYOP VDD VIN- VIN+ VOUT VSS
*.PININFO VDD:I VSS:I VIN-:I VIN+:I VOUT:I
xa1 net1 net1 VDD VDD JNWATR_PCH_4C1F2
xb1 net4 net1 VDD VDD JNWATR_PCH_4C1F2
xd VOUT net1 VDD VDD JNWATR_PCH_4C1F2
xd2 VOUT net3 VSS VSS JNWATR_NCH_4C1F2
xe net6 VDD net3 VSS JNWATR_NCH_2C1F2
xc2 net2 VIN- net4 net4 JNWATR_PCH_4C5F0
xc3 net2 net2 VSS VSS JNWATR_NCH_4C1F2
xb3 net3 net2 VSS VSS JNWATR_NCH_4C1F2
xb2 net3 VIN+ net4 net4 JNWATR_PCH_4C5F0
xa3 VSS net5 VSS JNWTR_RPPO16
xd1 net6 VOUT JNWTR_CAPX1
xa2 net5 net1 VSS JNWTR_RPPO2
.ends

* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sym # of pins=4
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sch
.subckt JNWATR_PCH_4C1F2 D G S B
*.PININFO D:B G:B S:B B:B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=3.2 nf=2 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C1F2.sym # of pins=4
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C1F2.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C1F2.sch
.subckt JNWATR_NCH_4C1F2 D G S B
*.PININFO D:B G:B S:B B:B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.22 W=3.2 nf=2 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_2C1F2.sym # of pins=4
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_2C1F2.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_2C1F2.sch
.subckt JNWATR_NCH_2C1F2 D G S B
*.PININFO D:B G:B S:B B:B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.22 W=1.92 nf=2 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym # of pins=4
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sch
.subckt JNWATR_PCH_4C5F0 D G S B
*.PININFO D:B G:B S:B B:B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=3.2 nf=2 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO16.sym # of pins=3
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO16.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO16.sch
.subckt JNWTR_RPPO16 N P B
*.PININFO P:B N:B B:B
XXA1 N P B JNWTR_RES16
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX1.sym # of pins=2
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sch
.subckt JNWTR_CAPX1 A B
*.PININFO A:B B:B
XC1 B A sky130_fd_pr__cap_mim_m3_1 W=5 L=5 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO2.sym # of pins=3
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO2.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO2.sch
.subckt JNWTR_RPPO2 N P B
*.PININFO P:B N:B B:B
XXA1 N P B JNWTR_RES2
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES16.sym # of pins=3
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RES16.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RES16.sch
.subckt JNWTR_RES16 N P B
*.PININFO N:B P:B B:B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 INT_3 INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_4 INT_4 INT_3 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_5 INT_5 INT_4 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_6 INT_6 INT_5 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_7 INT_7 INT_6 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_8 INT_8 INT_7 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_9 INT_9 INT_8 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_10 INT_10 INT_9 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_11 INT_11 INT_10 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_12 INT_12 INT_11 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_13 INT_13 INT_12 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_14 INT_14 INT_13 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_15 P INT_14 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES2.sym # of pins=3
** sym_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RES2.sym
** sch_path: /home/manu/pro/aicex/ip/jnw_gr01_sky130a/design/JNW_TR_SKY130A/JNWTR_RES2.sch
.subckt JNWTR_RES2 N P B
*.PININFO N:B P:B B:B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 P INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends

.end
